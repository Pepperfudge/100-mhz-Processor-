/**
 * UC Berkeley CS150
 * Fall 2014
 * List of ALU operations.
 */

`ifndef ALUOP
`define ALUOP

`define ALU_ADD     4'd0
`define ALU_SUB     4'd1
`define ALU_AND     4'd2
`define ALU_OR      4'd3
`define ALU_XOR     4'd4
`define ALU_SLT     4'd5
`define ALU_SLTU    4'd6
`define ALU_SLL     4'd7
`define ALU_SRA     4'd8
`define ALU_SRL     4'd9
`define ALU_COPY_B  4'd10
`define ALU_EQ      4'd11
`define ALU_NE      4'd12
`define ALU_GE      4'd13
`define ALU_GEU     4'd14
`define ALU_XXX     4'd15


`endif //ALUOP
