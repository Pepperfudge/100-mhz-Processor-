module asmtest(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h130f0000;
30'h00000001: inst = 32'h93030000;
30'h00000002: inst = 32'h93013000;
30'h00000003: inst = 32'h13024000;
30'h00000004: inst = 32'h93025000;
30'h00000005: inst = 32'h13036000;
30'h00000006: inst = 32'hb7000010;
30'h00000007: inst = 32'h93800002;
30'h00000008: inst = 32'h37b1ad1e;
30'h00000009: inst = 32'h1301f10e;
30'h0000000a: inst = 32'h37050010;
30'h0000000b: inst = 32'h23201500;
30'h0000000c: inst = 32'h23222500;
30'h0000000d: inst = 32'h83250500;
30'h0000000e: inst = 32'h03264500;
30'h0000000f: inst = 32'h930f1003;
30'h00000010: inst = 32'h93831300;
30'h00000011: inst = 32'h639eb05c;
30'h00000012: inst = 32'h930f2003;
30'h00000013: inst = 32'h93831300;
30'h00000014: inst = 32'h6318c15c;
30'h00000015: inst = 32'h930f3003;
30'h00000016: inst = 32'h93831300;
30'h00000017: inst = 32'h371a0000;
30'h00000018: inst = 32'h930a0040;
30'h00000019: inst = 32'h938a0a40;
30'h0000001a: inst = 32'h938a0a40;
30'h0000001b: inst = 32'h938a0a40;
30'h0000001c: inst = 32'h63984a5b;
30'h0000001d: inst = 32'h930f4003;
30'h0000001e: inst = 32'h93831300;
30'h0000001f: inst = 32'h930af04f;
30'h00000020: inst = 32'h136af04f;
30'h00000021: inst = 32'h639e4a59;
30'h00000022: inst = 32'h930f5003;
30'h00000023: inst = 32'h93831300;
30'h00000024: inst = 32'h170a0000;
30'h00000025: inst = 32'he70aca00;
30'h00000026: inst = 32'h6f00c062;
30'h00000027: inst = 32'h130a8a00;
30'h00000028: inst = 32'h63105a59;
30'h00000029: inst = 32'h930f6003;
30'h0000002a: inst = 32'h93831300;
30'h0000002b: inst = 32'h170a0000;
30'h0000002c: inst = 32'h135aca01;
30'h0000002d: inst = 32'h93021000;
30'h0000002e: inst = 32'h63944257;
30'h0000002f: inst = 32'h930f7003;
30'h00000030: inst = 32'h93831300;
30'h00000031: inst = 32'h130a1000;
30'h00000032: inst = 32'h930a2000;
30'h00000033: inst = 32'h130b2000;
30'h00000034: inst = 32'h630a5a5f;
30'h00000035: inst = 32'h63846a01;
30'h00000036: inst = 32'h6f008054;
30'h00000037: inst = 32'h930f8003;
30'h00000038: inst = 32'h93831300;
30'h00000039: inst = 32'h130a1000;
30'h0000003a: inst = 32'h930a2000;
30'h0000003b: inst = 32'hb7fbffff;
30'h0000003c: inst = 32'h63ca4a5d;
30'h0000003d: inst = 32'h63c87a5d;
30'h0000003e: inst = 32'h63c44b01;
30'h0000003f: inst = 32'h6f004052;
30'h00000040: inst = 32'h930f9003;
30'h00000041: inst = 32'h93831300;
30'h00000042: inst = 32'h130a1000;
30'h00000043: inst = 32'h930a2000;
30'h00000044: inst = 32'hb7fbffff;
30'h00000045: inst = 32'h63e84a5b;
30'h00000046: inst = 32'h63e64b5b;
30'h00000047: inst = 32'h63645a01;
30'h00000048: inst = 32'h6f000050;
30'h00000049: inst = 32'h930f1006;
30'h0000004a: inst = 32'h93831300;
30'h0000004b: inst = 32'h130a1000;
30'h0000004c: inst = 32'h930a2000;
30'h0000004d: inst = 32'hb7fbffff;
30'h0000004e: inst = 32'h63565a59;
30'h0000004f: inst = 32'h63d45b59;
30'h00000050: inst = 32'h63547a01;
30'h00000051: inst = 32'h6f00c04d;
30'h00000052: inst = 32'h930f2006;
30'h00000053: inst = 32'h93831300;
30'h00000054: inst = 32'h130a1000;
30'h00000055: inst = 32'h930a2000;
30'h00000056: inst = 32'hb7fbffff;
30'h00000057: inst = 32'h63747a57;
30'h00000058: inst = 32'h63725a57;
30'h00000059: inst = 32'h63705057;
30'h0000005a: inst = 32'h63f45b01;
30'h0000005b: inst = 32'h6f00404b;
30'h0000005c: inst = 32'h930f3006;
30'h0000005d: inst = 32'h93831300;
30'h0000005e: inst = 32'h130af00f;
30'h0000005f: inst = 32'h931a4a01;
30'h00000060: inst = 32'hb70bf00f;
30'h00000061: inst = 32'h639e5b49;
30'h00000062: inst = 32'h930f4006;
30'h00000063: inst = 32'h93831300;
30'h00000064: inst = 32'h37fcffff;
30'h00000065: inst = 32'h136cfcff;
30'h00000066: inst = 32'hb70b0080;
30'h00000067: inst = 32'h93dbfb41;
30'h00000068: inst = 32'h63107c49;
30'h00000069: inst = 32'h930f5006;
30'h0000006a: inst = 32'h93831300;
30'h0000006b: inst = 32'h37050010;
30'h0000006c: inst = 32'hb74a6587;
30'h0000006d: inst = 32'h93ea1a32;
30'h0000006e: inst = 32'h23205501;
30'h0000006f: inst = 32'h030b0500;
30'h00000070: inst = 32'h130c1002;
30'h00000071: inst = 32'h631e8b45;
30'h00000072: inst = 32'h030b1500;
30'h00000073: inst = 32'h130c3004;
30'h00000074: inst = 32'h63188b45;
30'h00000075: inst = 32'h030b2500;
30'h00000076: inst = 32'h130c5006;
30'h00000077: inst = 32'h63128b45;
30'h00000078: inst = 32'h030b3500;
30'h00000079: inst = 32'h370c0087;
30'h0000007a: inst = 32'h135c8c41;
30'h0000007b: inst = 32'h631a8b43;
30'h0000007c: inst = 32'h930f6006;
30'h0000007d: inst = 32'h93831300;
30'h0000007e: inst = 32'h37050010;
30'h0000007f: inst = 32'h370defcd;
30'h00000080: inst = 32'h135d0d01;
30'h00000081: inst = 32'h370aab89;
30'h00000082: inst = 32'hb3094d01;
30'h00000083: inst = 32'h23203501;
30'h00000084: inst = 32'h83270500;
30'h00000085: inst = 32'h030b0500;
30'h00000086: inst = 32'h370c00ef;
30'h00000087: inst = 32'h135c8c41;
30'h00000088: inst = 32'h63108b41;
30'h00000089: inst = 32'h030b1500;
30'h0000008a: inst = 32'h370c00cd;
30'h0000008b: inst = 32'h135c8c41;
30'h0000008c: inst = 32'h63188b3f;
30'h0000008d: inst = 32'h030b2500;
30'h0000008e: inst = 32'h370c00ab;
30'h0000008f: inst = 32'h135c8c41;
30'h00000090: inst = 32'h63108b3f;
30'h00000091: inst = 32'h832c0500;
30'h00000092: inst = 32'h030b3500;
30'h00000093: inst = 32'h370c0089;
30'h00000094: inst = 32'h135c8c41;
30'h00000095: inst = 32'h63168b3d;
30'h00000096: inst = 32'h930f7006;
30'h00000097: inst = 32'h93831300;
30'h00000098: inst = 32'h37050010;
30'h00000099: inst = 32'h370defcd;
30'h0000009a: inst = 32'h135d0d01;
30'h0000009b: inst = 32'h370aab89;
30'h0000009c: inst = 32'hb3094d01;
30'h0000009d: inst = 32'h23203501;
30'h0000009e: inst = 32'h83270500;
30'h0000009f: inst = 32'h031b0500;
30'h000000a0: inst = 32'h370cefcd;
30'h000000a1: inst = 32'h135c0c41;
30'h000000a2: inst = 32'h631c8b39;
30'h000000a3: inst = 32'h031b2500;
30'h000000a4: inst = 32'h370cab89;
30'h000000a5: inst = 32'h135c0c41;
30'h000000a6: inst = 32'h63148b39;
30'h000000a7: inst = 32'h930f8006;
30'h000000a8: inst = 32'h93831300;
30'h000000a9: inst = 32'h37050010;
30'h000000aa: inst = 32'h370d2143;
30'h000000ab: inst = 32'h135d0d01;
30'h000000ac: inst = 32'h370a6587;
30'h000000ad: inst = 32'hb3094d01;
30'h000000ae: inst = 32'h23203501;
30'h000000af: inst = 32'h83270500;
30'h000000b0: inst = 32'h031b0500;
30'h000000b1: inst = 32'h370c2143;
30'h000000b2: inst = 32'h135c0c41;
30'h000000b3: inst = 32'h631a8b35;
30'h000000b4: inst = 32'h031b2500;
30'h000000b5: inst = 32'h370c6587;
30'h000000b6: inst = 32'h135c0c41;
30'h000000b7: inst = 32'h63128b35;
30'h000000b8: inst = 32'h930f9006;
30'h000000b9: inst = 32'h93831300;
30'h000000ba: inst = 32'h37050010;
30'h000000bb: inst = 32'h370d2143;
30'h000000bc: inst = 32'h135d0d01;
30'h000000bd: inst = 32'h370a6587;
30'h000000be: inst = 32'hb3094d01;
30'h000000bf: inst = 32'h23203501;
30'h000000c0: inst = 32'h83270500;
30'h000000c1: inst = 32'h639e3731;
30'h000000c2: inst = 32'h930fa006;
30'h000000c3: inst = 32'h93831300;
30'h000000c4: inst = 32'h37050010;
30'h000000c5: inst = 32'hb74a6587;
30'h000000c6: inst = 32'h93ea1a32;
30'h000000c7: inst = 32'h23205501;
30'h000000c8: inst = 32'h034b0500;
30'h000000c9: inst = 32'h130c1002;
30'h000000ca: inst = 32'h631c8b2f;
30'h000000cb: inst = 32'h034b1500;
30'h000000cc: inst = 32'h130c3004;
30'h000000cd: inst = 32'h63168b2f;
30'h000000ce: inst = 32'h034b2500;
30'h000000cf: inst = 32'h130c5006;
30'h000000d0: inst = 32'h63108b2f;
30'h000000d1: inst = 32'h034b3500;
30'h000000d2: inst = 32'h370c0087;
30'h000000d3: inst = 32'h135c8c01;
30'h000000d4: inst = 32'h63188b2d;
30'h000000d5: inst = 32'h930fb006;
30'h000000d6: inst = 32'h93831300;
30'h000000d7: inst = 32'h37050010;
30'h000000d8: inst = 32'h370defcd;
30'h000000d9: inst = 32'h135d0d01;
30'h000000da: inst = 32'h370aab89;
30'h000000db: inst = 32'hb3094d01;
30'h000000dc: inst = 32'h23203501;
30'h000000dd: inst = 32'h83270500;
30'h000000de: inst = 32'h034b0500;
30'h000000df: inst = 32'h370c00ef;
30'h000000e0: inst = 32'h135c8c01;
30'h000000e1: inst = 32'h631e8b29;
30'h000000e2: inst = 32'h034b1500;
30'h000000e3: inst = 32'h370c00cd;
30'h000000e4: inst = 32'h135c8c01;
30'h000000e5: inst = 32'h63168b29;
30'h000000e6: inst = 32'h034b2500;
30'h000000e7: inst = 32'h370c00ab;
30'h000000e8: inst = 32'h135c8c01;
30'h000000e9: inst = 32'h631e8b27;
30'h000000ea: inst = 32'h034b3500;
30'h000000eb: inst = 32'h370c0089;
30'h000000ec: inst = 32'h135c8c01;
30'h000000ed: inst = 32'h63168b27;
30'h000000ee: inst = 32'h930fc006;
30'h000000ef: inst = 32'h93831300;
30'h000000f0: inst = 32'h37050010;
30'h000000f1: inst = 32'h370defcd;
30'h000000f2: inst = 32'h135d0d01;
30'h000000f3: inst = 32'h370aab89;
30'h000000f4: inst = 32'hb3094d01;
30'h000000f5: inst = 32'h23203501;
30'h000000f6: inst = 32'h83270500;
30'h000000f7: inst = 32'h035b0500;
30'h000000f8: inst = 32'h370cefcd;
30'h000000f9: inst = 32'h135c0c01;
30'h000000fa: inst = 32'h631c8b23;
30'h000000fb: inst = 32'h035b2500;
30'h000000fc: inst = 32'h370cab89;
30'h000000fd: inst = 32'h135c0c01;
30'h000000fe: inst = 32'h63148b23;
30'h000000ff: inst = 32'h930fd006;
30'h00000100: inst = 32'h93831300;
30'h00000101: inst = 32'h37050010;
30'h00000102: inst = 32'h370d2143;
30'h00000103: inst = 32'h135d0d01;
30'h00000104: inst = 32'h370a6587;
30'h00000105: inst = 32'hb3094d01;
30'h00000106: inst = 32'h23203501;
30'h00000107: inst = 32'h83270500;
30'h00000108: inst = 32'h035b0500;
30'h00000109: inst = 32'h370c2143;
30'h0000010a: inst = 32'h135c0c01;
30'h0000010b: inst = 32'h631a8b1f;
30'h0000010c: inst = 32'h035b2500;
30'h0000010d: inst = 32'h370c6587;
30'h0000010e: inst = 32'h135c0c01;
30'h0000010f: inst = 32'h63128b1f;
30'h00000110: inst = 32'h930fe006;
30'h00000111: inst = 32'h93831300;
30'h00000112: inst = 32'h37050010;
30'h00000113: inst = 32'h370d2143;
30'h00000114: inst = 32'h135d0d01;
30'h00000115: inst = 32'h370a6587;
30'h00000116: inst = 32'hb3094d01;
30'h00000117: inst = 32'h23200500;
30'h00000118: inst = 32'h23003501;
30'h00000119: inst = 32'h370c0021;
30'h0000011a: inst = 32'h135c8c01;
30'h0000011b: inst = 32'h032b0500;
30'h0000011c: inst = 32'h63188b1b;
30'h0000011d: inst = 32'ha3003501;
30'h0000011e: inst = 32'h370c2121;
30'h0000011f: inst = 32'h135c0c01;
30'h00000120: inst = 32'h032b0500;
30'h00000121: inst = 32'h631e8b19;
30'h00000122: inst = 32'h23200500;
30'h00000123: inst = 32'h23013501;
30'h00000124: inst = 32'h370c2100;
30'h00000125: inst = 32'h032b0500;
30'h00000126: inst = 32'h63148b19;
30'h00000127: inst = 32'ha3013501;
30'h00000128: inst = 32'h370c2121;
30'h00000129: inst = 32'h032b0500;
30'h0000012a: inst = 32'h631c8b17;
30'h0000012b: inst = 32'h930fe006;
30'h0000012c: inst = 32'h93831300;
30'h0000012d: inst = 32'h37050010;
30'h0000012e: inst = 32'h370d2143;
30'h0000012f: inst = 32'h135d0d01;
30'h00000130: inst = 32'h370a6587;
30'h00000131: inst = 32'hb3094d01;
30'h00000132: inst = 32'h23200500;
30'h00000133: inst = 32'h23003501;
30'h00000134: inst = 32'h370c0021;
30'h00000135: inst = 32'h135c8c01;
30'h00000136: inst = 32'h032b0500;
30'h00000137: inst = 32'h63128b15;
30'h00000138: inst = 32'ha3003501;
30'h00000139: inst = 32'h370c2121;
30'h0000013a: inst = 32'h135c0c01;
30'h0000013b: inst = 32'h032b0500;
30'h0000013c: inst = 32'h63188b13;
30'h0000013d: inst = 32'h23200500;
30'h0000013e: inst = 32'h23013501;
30'h0000013f: inst = 32'h370c2100;
30'h00000140: inst = 32'h032b0500;
30'h00000141: inst = 32'h631e8b11;
30'h00000142: inst = 32'ha3013501;
30'h00000143: inst = 32'h370c2121;
30'h00000144: inst = 32'h032b0500;
30'h00000145: inst = 32'h63168b11;
30'h00000146: inst = 32'h930fc006;
30'h00000147: inst = 32'h93831300;
30'h00000148: inst = 32'h370d2143;
30'h00000149: inst = 32'h135d0d01;
30'h0000014a: inst = 32'h370a6587;
30'h0000014b: inst = 32'hb3094d01;
30'h0000014c: inst = 32'h23223501;
30'h0000014d: inst = 32'h032b4500;
30'h0000014e: inst = 32'h6394690f;
30'h0000014f: inst = 32'h930ff006;
30'h00000150: inst = 32'h93831300;
30'h00000151: inst = 32'h37050010;
30'h00000152: inst = 32'h370d2143;
30'h00000153: inst = 32'h135d0d01;
30'h00000154: inst = 32'h370a6587;
30'h00000155: inst = 32'hb3094d01;
30'h00000156: inst = 32'h23203501;
30'h00000157: inst = 32'h370d3412;
30'h00000158: inst = 32'h135d0d01;
30'h00000159: inst = 32'h2310a501;
30'h0000015a: inst = 32'h032b0500;
30'h0000015b: inst = 32'h370d3412;
30'h0000015c: inst = 32'h135d0d01;
30'h0000015d: inst = 32'h370a6587;
30'h0000015e: inst = 32'h330c4d01;
30'h0000015f: inst = 32'h63128b0b;
30'h00000160: inst = 32'h370d2143;
30'h00000161: inst = 32'h135d0d01;
30'h00000162: inst = 32'h2311a501;
30'h00000163: inst = 32'h032b0500;
30'h00000164: inst = 32'hb70c3412;
30'h00000165: inst = 32'h93dc0c01;
30'h00000166: inst = 32'h370a2143;
30'h00000167: inst = 32'h338c4c01;
30'h00000168: inst = 32'h63108b09;
30'h00000169: inst = 32'h930f0007;
30'h0000016a: inst = 32'h93831300;
30'h0000016b: inst = 32'h37050010;
30'h0000016c: inst = 32'h93054500;
30'h0000016d: inst = 32'h130d5000;
30'h0000016e: inst = 32'h23aea5ff;
30'h0000016f: inst = 32'h83220500;
30'h00000170: inst = 32'h6390a207;
30'h00000171: inst = 32'h930f1007;
30'h00000172: inst = 32'h93831300;
30'h00000173: inst = 32'hef00c000;
30'h00000174: inst = 32'h03a40500;
30'h00000175: inst = 32'h63166404;
30'h00000176: inst = 32'h13036000;
30'h00000177: inst = 32'hb7050010;
30'h00000178: inst = 32'h13050040;
30'h00000179: inst = 32'h13158500;
30'h0000017a: inst = 32'hb305b500;
30'h0000017b: inst = 32'h23a06500;
30'h0000017c: inst = 32'he7800000;
30'h0000017d: inst = 32'h930f2007;
30'h0000017e: inst = 32'h93831300;
30'h0000017f: inst = 32'h13012000;
30'h00000180: inst = 32'h330a0000;
30'h00000181: inst = 32'h63040000;
30'h00000182: inst = 32'h130aaa00;
30'h00000183: inst = 32'h33000000;
30'h00000184: inst = 32'h33000000;
30'h00000185: inst = 32'h130a2a00;
30'h00000186: inst = 32'h63144101;
30'h00000187: inst = 32'h6f00c00e;
30'h00000188: inst = 32'h13026004;
30'h00000189: inst = 32'hef008017;
30'h0000018a: inst = 32'h13021004;
30'h0000018b: inst = 32'hef000017;
30'h0000018c: inst = 32'h13029004;
30'h0000018d: inst = 32'hef008016;
30'h0000018e: inst = 32'h1302c004;
30'h0000018f: inst = 32'hef000016;
30'h00000190: inst = 32'h13026004;
30'h00000191: inst = 32'hef008015;
30'h00000192: inst = 32'h13021004;
30'h00000193: inst = 32'hef000015;
30'h00000194: inst = 32'h13029004;
30'h00000195: inst = 32'hef008014;
30'h00000196: inst = 32'h1302c004;
30'h00000197: inst = 32'hef000014;
30'h00000198: inst = 32'h13026004;
30'h00000199: inst = 32'hef008013;
30'h0000019a: inst = 32'h13021004;
30'h0000019b: inst = 32'hef000013;
30'h0000019c: inst = 32'h13029004;
30'h0000019d: inst = 32'hef008012;
30'h0000019e: inst = 32'h1302c004;
30'h0000019f: inst = 32'hef000012;
30'h000001a0: inst = 32'h13026004;
30'h000001a1: inst = 32'hef008011;
30'h000001a2: inst = 32'h13021004;
30'h000001a3: inst = 32'hef000011;
30'h000001a4: inst = 32'h13029004;
30'h000001a5: inst = 32'hef008010;
30'h000001a6: inst = 32'h1302c004;
30'h000001a7: inst = 32'hef000010;
30'h000001a8: inst = 32'h1302a003;
30'h000001a9: inst = 32'hef00800f;
30'h000001aa: inst = 32'h13020002;
30'h000001ab: inst = 32'hef00000f;
30'h000001ac: inst = 32'h3302f001;
30'h000001ad: inst = 32'hef00800e;
30'h000001ae: inst = 32'h1302a000;
30'h000001af: inst = 32'hef00000e;
30'h000001b0: inst = 32'h6f00400d;
30'h000001b1: inst = 32'h13026004;
30'h000001b2: inst = 32'hef00400d;
30'h000001b3: inst = 32'h1302c004;
30'h000001b4: inst = 32'hef00c00c;
30'h000001b5: inst = 32'h13021004;
30'h000001b6: inst = 32'hef00400c;
30'h000001b7: inst = 32'h13027004;
30'h000001b8: inst = 32'hef00c00b;
30'h000001b9: inst = 32'h1302a003;
30'h000001ba: inst = 32'hef00400b;
30'h000001bb: inst = 32'h13020002;
30'h000001bc: inst = 32'hef00c00a;
30'h000001bd: inst = 32'h3302f001;
30'h000001be: inst = 32'hef00400a;
30'h000001bf: inst = 32'h1302a000;
30'h000001c0: inst = 32'hef00c009;
30'h000001c1: inst = 32'h6f000009;
30'h000001c2: inst = 32'h13020005;
30'h000001c3: inst = 32'hef000009;
30'h000001c4: inst = 32'h13021004;
30'h000001c5: inst = 32'hef008008;
30'h000001c6: inst = 32'h13023005;
30'h000001c7: inst = 32'hef000008;
30'h000001c8: inst = 32'h13023005;
30'h000001c9: inst = 32'hef008007;
30'h000001ca: inst = 32'h13020005;
30'h000001cb: inst = 32'hef000007;
30'h000001cc: inst = 32'h13021004;
30'h000001cd: inst = 32'hef008006;
30'h000001ce: inst = 32'h13023005;
30'h000001cf: inst = 32'hef000006;
30'h000001d0: inst = 32'h13023005;
30'h000001d1: inst = 32'hef008005;
30'h000001d2: inst = 32'h13020005;
30'h000001d3: inst = 32'hef000005;
30'h000001d4: inst = 32'h13021004;
30'h000001d5: inst = 32'hef008004;
30'h000001d6: inst = 32'h13023005;
30'h000001d7: inst = 32'hef000004;
30'h000001d8: inst = 32'h13023005;
30'h000001d9: inst = 32'hef008003;
30'h000001da: inst = 32'h13020005;
30'h000001db: inst = 32'hef000003;
30'h000001dc: inst = 32'h13021004;
30'h000001dd: inst = 32'hef008002;
30'h000001de: inst = 32'h13023005;
30'h000001df: inst = 32'hef000002;
30'h000001e0: inst = 32'h13023005;
30'h000001e1: inst = 32'hef008001;
30'h000001e2: inst = 32'h1302a000;
30'h000001e3: inst = 32'hef000001;
30'h000001e4: inst = 32'h6f004000;
30'h000001e5: inst = 32'h130f1000;
30'h000001e6: inst = 32'h6ff0dfff;
30'h000001e7: inst = 32'h37010080;
30'h000001e8: inst = 32'h83210100;
30'h000001e9: inst = 32'h93f11100;
30'h000001ea: inst = 32'he38a01fe;
30'h000001eb: inst = 32'h23244100;
30'h000001ec: inst = 32'h67800000;
default:      inst = 32'h00000000;
endcase
end
endmodule
