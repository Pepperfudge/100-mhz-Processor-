module asmtest(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h93037000;
30'h00000001: inst = 32'h93001000;
30'h00000002: inst = 32'h13012000;
30'h00000003: inst = 32'h33841300;
30'h00000004: inst = 32'hb3041400;
30'h00000005: inst = 32'h33859000;
30'h00000006: inst = 32'hb70f0080;
30'h00000007: inst = 32'h938f1f00;
30'h00000008: inst = 32'h970f0080;
30'h00000009: inst = 32'hb38f0f00;
30'h0000000a: inst = 32'h638c7300;
30'h0000000b: inst = 32'hb70f0080;
30'h0000000c: inst = 32'h13000000;
30'h0000000d: inst = 32'h13000000;
30'h0000000e: inst = 32'h13000000;
30'h0000000f: inst = 32'h13000000;
30'h00000010: inst = 32'h93051500;
30'h00000011: inst = 32'hef008000;
30'h00000012: inst = 32'h33000000;
30'h00000013: inst = 32'h93800000;
30'h00000014: inst = 32'h93001000;
30'h00000015: inst = 32'h37050010;
30'h00000016: inst = 32'h23201500;
30'h00000017: inst = 32'h23222500;
30'h00000018: inst = 32'h83250500;
30'h00000019: inst = 32'h03264500;
30'h0000001a: inst = 32'h13010600;
30'h0000001b: inst = 32'h93800500;
default:      inst = 32'h00000000;
endcase
end
endmodule
