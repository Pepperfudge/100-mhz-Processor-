module asmtest(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h37050030;
30'h00000001: inst = 32'hb7100000;
30'h00000002: inst = 32'h938030f1;
30'h00000003: inst = 32'h3705ff3f;
30'h00000004: inst = 32'h23201500;
30'h00000005: inst = 32'h93003039;
30'h00000006: inst = 32'h3705ff3f;
30'h00000007: inst = 32'h13054500;
30'h00000008: inst = 32'h23201500;
30'h00000009: inst = 32'hb7003000;
30'h0000000a: inst = 32'h93803019;
30'h0000000b: inst = 32'h3705ff3f;
30'h0000000c: inst = 32'h13058500;
30'h0000000d: inst = 32'h23201500;
30'h0000000e: inst = 32'hb7004000;
30'h0000000f: inst = 32'h93803021;
30'h00000010: inst = 32'h3705ff3f;
30'h00000011: inst = 32'h1305c500;
30'h00000012: inst = 32'h23201500;
30'h00000013: inst = 32'hb7005000;
30'h00000014: inst = 32'h93803029;
30'h00000015: inst = 32'h3705ff3f;
30'h00000016: inst = 32'h13050501;
30'h00000017: inst = 32'h23201500;
30'h00000018: inst = 32'hb7006000;
30'h00000019: inst = 32'h93803031;
30'h0000001a: inst = 32'h3705ff3f;
30'h0000001b: inst = 32'h13054501;
30'h0000001c: inst = 32'h23201500;
30'h0000001d: inst = 32'hb7000010;
30'h0000001e: inst = 32'h9380700b;
30'h0000001f: inst = 32'h3705ff3f;
30'h00000020: inst = 32'h13058501;
30'h00000021: inst = 32'h23201500;
30'h00000022: inst = 32'hb7800002;
30'h00000023: inst = 32'h93803009;
30'h00000024: inst = 32'h3705ff3f;
30'h00000025: inst = 32'h1305c501;
30'h00000026: inst = 32'h23201500;
30'h00000027: inst = 32'hb7b0ad1e;
30'h00000028: inst = 32'h93807013;
30'h00000029: inst = 32'h3705ff3f;
30'h0000002a: inst = 32'h13050502;
30'h0000002b: inst = 32'h23201500;
30'h0000002c: inst = 32'hb700f10e;
30'h0000002d: inst = 32'h93803011;
30'h0000002e: inst = 32'h3705ff3f;
30'h0000002f: inst = 32'h13054502;
30'h00000030: inst = 32'h23201500;
30'h00000031: inst = 32'hb7000010;
30'h00000032: inst = 32'h93807053;
30'h00000033: inst = 32'h3705ff3f;
30'h00000034: inst = 32'h13058502;
30'h00000035: inst = 32'h23201500;
30'h00000036: inst = 32'hb7201500;
30'h00000037: inst = 32'h93803002;
30'h00000038: inst = 32'h3705ff3f;
30'h00000039: inst = 32'h1305c502;
30'h0000003a: inst = 32'h23201500;
30'h0000003b: inst = 32'hb7202500;
30'h0000003c: inst = 32'h93803022;
30'h0000003d: inst = 32'h3705ff3f;
30'h0000003e: inst = 32'h13050503;
30'h0000003f: inst = 32'h23201500;
30'h00000040: inst = 32'hb7200500;
30'h00000041: inst = 32'h93803058;
30'h00000042: inst = 32'h3705ff3f;
30'h00000043: inst = 32'h13054503;
30'h00000044: inst = 32'h23201500;
30'h00000045: inst = 32'hb7204500;
30'h00000046: inst = 32'h93803060;
30'h00000047: inst = 32'h3705ff3f;
30'h00000048: inst = 32'h13058503;
30'h00000049: inst = 32'h23201500;
30'h0000004a: inst = 32'hb7101003;
30'h0000004b: inst = 32'h938030f9;
30'h0000004c: inst = 32'h3705ff3f;
30'h0000004d: inst = 32'h1305c503;
30'h0000004e: inst = 32'h23201500;
30'h0000004f: inst = 32'hb7801300;
30'h00000050: inst = 32'h93803039;
30'h00000051: inst = 32'h3705ff3f;
30'h00000052: inst = 32'h13050504;
30'h00000053: inst = 32'h23201500;
30'h00000054: inst = 32'hb7a0b05c;
30'h00000055: inst = 32'h938030e6;
30'h00000056: inst = 32'h3705ff3f;
30'h00000057: inst = 32'h13054504;
30'h00000058: inst = 32'h23201500;
30'h00000059: inst = 32'hb7102003;
30'h0000005a: inst = 32'h938030f9;
30'h0000005b: inst = 32'h3705ff3f;
30'h0000005c: inst = 32'h13058504;
30'h0000005d: inst = 32'h23201500;
30'h0000005e: inst = 32'hb7801300;
30'h0000005f: inst = 32'h93803039;
30'h00000060: inst = 32'h3705ff3f;
30'h00000061: inst = 32'h1305c504;
30'h00000062: inst = 32'h23201500;
30'h00000063: inst = 32'hb720c15c;
30'h00000064: inst = 32'h93803086;
30'h00000065: inst = 32'h3705ff3f;
30'h00000066: inst = 32'h13050505;
30'h00000067: inst = 32'h23201500;
30'h00000068: inst = 32'hb7103003;
30'h00000069: inst = 32'h938030f9;
30'h0000006a: inst = 32'h3705ff3f;
30'h0000006b: inst = 32'h13054505;
30'h0000006c: inst = 32'h23201500;
30'h0000006d: inst = 32'hb7801300;
30'h0000006e: inst = 32'h93803039;
30'h0000006f: inst = 32'h3705ff3f;
30'h00000070: inst = 32'h13058505;
30'h00000071: inst = 32'h23201500;
30'h00000072: inst = 32'hb7200000;
30'h00000073: inst = 32'h938070a3;
30'h00000074: inst = 32'h3705ff3f;
30'h00000075: inst = 32'h1305c505;
30'h00000076: inst = 32'h23201500;
30'h00000077: inst = 32'hb7100040;
30'h00000078: inst = 32'h938030a9;
30'h00000079: inst = 32'h3705ff3f;
30'h0000007a: inst = 32'h13050506;
30'h0000007b: inst = 32'h23201500;
30'h0000007c: inst = 32'hb7900a40;
30'h0000007d: inst = 32'h938030a9;
30'h0000007e: inst = 32'h3705ff3f;
30'h0000007f: inst = 32'h13054506;
30'h00000080: inst = 32'h23201500;
30'h00000081: inst = 32'hb7900a40;
30'h00000082: inst = 32'h938030a9;
30'h00000083: inst = 32'h3705ff3f;
30'h00000084: inst = 32'h13058506;
30'h00000085: inst = 32'h23201500;
30'h00000086: inst = 32'hb7900a40;
30'h00000087: inst = 32'h938030a9;
30'h00000088: inst = 32'h3705ff3f;
30'h00000089: inst = 32'h1305c506;
30'h0000008a: inst = 32'h23201500;
30'h0000008b: inst = 32'hb7a04a5b;
30'h0000008c: inst = 32'h93803086;
30'h0000008d: inst = 32'h3705ff3f;
30'h0000008e: inst = 32'h13050507;
30'h0000008f: inst = 32'h23201500;
30'h00000090: inst = 32'hb7104003;
30'h00000091: inst = 32'h938030f9;
30'h00000092: inst = 32'h3705ff3f;
30'h00000093: inst = 32'h13054507;
30'h00000094: inst = 32'h23201500;
30'h00000095: inst = 32'hb7801300;
30'h00000096: inst = 32'h93803039;
30'h00000097: inst = 32'h3705ff3f;
30'h00000098: inst = 32'h13058507;
30'h00000099: inst = 32'h23201500;
30'h0000009a: inst = 32'hb710f04f;
30'h0000009b: inst = 32'h938030a9;
30'h0000009c: inst = 32'h3705ff3f;
30'h0000009d: inst = 32'h1305c507;
30'h0000009e: inst = 32'h23201500;
30'h0000009f: inst = 32'hb770f04f;
30'h000000a0: inst = 32'h938030a1;
30'h000000a1: inst = 32'h3705ff3f;
30'h000000a2: inst = 32'h13050508;
30'h000000a3: inst = 32'h23201500;
30'h000000a4: inst = 32'hb7a04a59;
30'h000000a5: inst = 32'h938030e6;
30'h000000a6: inst = 32'h3705ff3f;
30'h000000a7: inst = 32'h13054508;
30'h000000a8: inst = 32'h23201500;
30'h000000a9: inst = 32'hb7105003;
30'h000000aa: inst = 32'h938030f9;
30'h000000ab: inst = 32'h3705ff3f;
30'h000000ac: inst = 32'h13058508;
30'h000000ad: inst = 32'h23201500;
30'h000000ae: inst = 32'hb7801300;
30'h000000af: inst = 32'h93803039;
30'h000000b0: inst = 32'h3705ff3f;
30'h000000b1: inst = 32'h1305c508;
30'h000000b2: inst = 32'h23201500;
30'h000000b3: inst = 32'hb7100000;
30'h000000b4: inst = 32'h938070a1;
30'h000000b5: inst = 32'h3705ff3f;
30'h000000b6: inst = 32'h13050509;
30'h000000b7: inst = 32'h23201500;
30'h000000b8: inst = 32'hb710ca00;
30'h000000b9: inst = 32'h938070ae;
30'h000000ba: inst = 32'h3705ff3f;
30'h000000bb: inst = 32'h13054509;
30'h000000bc: inst = 32'h23201500;
30'h000000bd: inst = 32'hb700c062;
30'h000000be: inst = 32'h9380f006;
30'h000000bf: inst = 32'h3705ff3f;
30'h000000c0: inst = 32'h13058509;
30'h000000c1: inst = 32'h23201500;
30'h000000c2: inst = 32'hb7108a00;
30'h000000c3: inst = 32'h938030a1;
30'h000000c4: inst = 32'h3705ff3f;
30'h000000c5: inst = 32'h1305c509;
30'h000000c6: inst = 32'h23201500;
30'h000000c7: inst = 32'hb7105a59;
30'h000000c8: inst = 32'h93803006;
30'h000000c9: inst = 32'h3705ff3f;
30'h000000ca: inst = 32'h1305050a;
30'h000000cb: inst = 32'h23201500;
30'h000000cc: inst = 32'hb7106003;
30'h000000cd: inst = 32'h938030f9;
30'h000000ce: inst = 32'h3705ff3f;
30'h000000cf: inst = 32'h1305450a;
30'h000000d0: inst = 32'h23201500;
30'h000000d1: inst = 32'hb7801300;
30'h000000d2: inst = 32'h93803039;
30'h000000d3: inst = 32'h3705ff3f;
30'h000000d4: inst = 32'h1305850a;
30'h000000d5: inst = 32'h23201500;
30'h000000d6: inst = 32'hb7100000;
30'h000000d7: inst = 32'h938070a1;
30'h000000d8: inst = 32'h3705ff3f;
30'h000000d9: inst = 32'h1305c50a;
30'h000000da: inst = 32'h23201500;
30'h000000db: inst = 32'hb760ca01;
30'h000000dc: inst = 32'h938030a1;
30'h000000dd: inst = 32'h3705ff3f;
30'h000000de: inst = 32'h1305050b;
30'h000000df: inst = 32'h23201500;
30'h000000e0: inst = 32'hb7001000;
30'h000000e1: inst = 32'h93803029;
30'h000000e2: inst = 32'h3705ff3f;
30'h000000e3: inst = 32'h1305450b;
30'h000000e4: inst = 32'h23201500;
30'h000000e5: inst = 32'hb7904257;
30'h000000e6: inst = 32'h93803046;
30'h000000e7: inst = 32'h3705ff3f;
30'h000000e8: inst = 32'h1305850b;
30'h000000e9: inst = 32'h23201500;
30'h000000ea: inst = 32'hb7107003;
30'h000000eb: inst = 32'h938030f9;
30'h000000ec: inst = 32'h3705ff3f;
30'h000000ed: inst = 32'h1305c50b;
30'h000000ee: inst = 32'h23201500;
30'h000000ef: inst = 32'hb7801300;
30'h000000f0: inst = 32'h93803039;
30'h000000f1: inst = 32'h3705ff3f;
30'h000000f2: inst = 32'h1305050c;
30'h000000f3: inst = 32'h23201500;
30'h000000f4: inst = 32'hb7101000;
30'h000000f5: inst = 32'h938030a1;
30'h000000f6: inst = 32'h3705ff3f;
30'h000000f7: inst = 32'h1305450c;
30'h000000f8: inst = 32'h23201500;
30'h000000f9: inst = 32'hb7102000;
30'h000000fa: inst = 32'h938030a9;
30'h000000fb: inst = 32'h3705ff3f;
30'h000000fc: inst = 32'h1305850c;
30'h000000fd: inst = 32'h23201500;
30'h000000fe: inst = 32'hb7102000;
30'h000000ff: inst = 32'h938030b1;
30'h00000100: inst = 32'h3705ff3f;
30'h00000101: inst = 32'h1305c50c;
30'h00000102: inst = 32'h23201500;
30'h00000103: inst = 32'hb7105a5f;
30'h00000104: inst = 32'h938030a6;
30'h00000105: inst = 32'h3705ff3f;
30'h00000106: inst = 32'h1305050d;
30'h00000107: inst = 32'h23201500;
30'h00000108: inst = 32'hb7806a01;
30'h00000109: inst = 32'h93803046;
30'h0000010a: inst = 32'h3705ff3f;
30'h0000010b: inst = 32'h1305450d;
30'h0000010c: inst = 32'h23201500;
30'h0000010d: inst = 32'hb7008054;
30'h0000010e: inst = 32'h9380f006;
30'h0000010f: inst = 32'h3705ff3f;
30'h00000110: inst = 32'h1305850d;
30'h00000111: inst = 32'h23201500;
30'h00000112: inst = 32'hb7108003;
30'h00000113: inst = 32'h938030f9;
30'h00000114: inst = 32'h3705ff3f;
30'h00000115: inst = 32'h1305c50d;
30'h00000116: inst = 32'h23201500;
30'h00000117: inst = 32'hb7801300;
30'h00000118: inst = 32'h93803039;
30'h00000119: inst = 32'h3705ff3f;
30'h0000011a: inst = 32'h1305050e;
30'h0000011b: inst = 32'h23201500;
30'h0000011c: inst = 32'hb7101000;
30'h0000011d: inst = 32'h938030a1;
30'h0000011e: inst = 32'h3705ff3f;
30'h0000011f: inst = 32'h1305450e;
30'h00000120: inst = 32'h23201500;
30'h00000121: inst = 32'hb7102000;
30'h00000122: inst = 32'h938030a9;
30'h00000123: inst = 32'h3705ff3f;
30'h00000124: inst = 32'h1305850e;
30'h00000125: inst = 32'h23201500;
30'h00000126: inst = 32'h930070bb;
30'h00000127: inst = 32'h3705ff3f;
30'h00000128: inst = 32'h1305c50e;
30'h00000129: inst = 32'h23201500;
30'h0000012a: inst = 32'hb7d04a5d;
30'h0000012b: inst = 32'h938030a6;
30'h0000012c: inst = 32'h3705ff3f;
30'h0000012d: inst = 32'h1305050f;
30'h0000012e: inst = 32'h23201500;
30'h0000012f: inst = 32'hb7d07a5d;
30'h00000130: inst = 32'h93803086;
30'h00000131: inst = 32'h3705ff3f;
30'h00000132: inst = 32'h1305450f;
30'h00000133: inst = 32'h23201500;
30'h00000134: inst = 32'hb7c04b01;
30'h00000135: inst = 32'h93803046;
30'h00000136: inst = 32'h3705ff3f;
30'h00000137: inst = 32'h1305850f;
30'h00000138: inst = 32'h23201500;
30'h00000139: inst = 32'hb7004052;
30'h0000013a: inst = 32'h9380f006;
30'h0000013b: inst = 32'h3705ff3f;
30'h0000013c: inst = 32'h1305c50f;
30'h0000013d: inst = 32'h23201500;
30'h0000013e: inst = 32'hb7109003;
30'h0000013f: inst = 32'h938030f9;
30'h00000140: inst = 32'h3705ff3f;
30'h00000141: inst = 32'h13050510;
30'h00000142: inst = 32'h23201500;
30'h00000143: inst = 32'hb7801300;
30'h00000144: inst = 32'h93803039;
30'h00000145: inst = 32'h3705ff3f;
30'h00000146: inst = 32'h13054510;
30'h00000147: inst = 32'h23201500;
30'h00000148: inst = 32'hb7101000;
30'h00000149: inst = 32'h938030a1;
30'h0000014a: inst = 32'h3705ff3f;
30'h0000014b: inst = 32'h13058510;
30'h0000014c: inst = 32'h23201500;
30'h0000014d: inst = 32'hb7102000;
30'h0000014e: inst = 32'h938030a9;
30'h0000014f: inst = 32'h3705ff3f;
30'h00000150: inst = 32'h1305c510;
30'h00000151: inst = 32'h23201500;
30'h00000152: inst = 32'h930070bb;
30'h00000153: inst = 32'h3705ff3f;
30'h00000154: inst = 32'h13050511;
30'h00000155: inst = 32'h23201500;
30'h00000156: inst = 32'hb7f04a5b;
30'h00000157: inst = 32'h93803086;
30'h00000158: inst = 32'h3705ff3f;
30'h00000159: inst = 32'h13054511;
30'h0000015a: inst = 32'h23201500;
30'h0000015b: inst = 32'hb7e04b5b;
30'h0000015c: inst = 32'h93803066;
30'h0000015d: inst = 32'h3705ff3f;
30'h0000015e: inst = 32'h13058511;
30'h0000015f: inst = 32'h23201500;
30'h00000160: inst = 32'hb7605a01;
30'h00000161: inst = 32'h93803046;
30'h00000162: inst = 32'h3705ff3f;
30'h00000163: inst = 32'h1305c511;
30'h00000164: inst = 32'h23201500;
30'h00000165: inst = 32'hb7000050;
30'h00000166: inst = 32'h9380f006;
30'h00000167: inst = 32'h3705ff3f;
30'h00000168: inst = 32'h13050512;
30'h00000169: inst = 32'h23201500;
30'h0000016a: inst = 32'hb7101006;
30'h0000016b: inst = 32'h938030f9;
30'h0000016c: inst = 32'h3705ff3f;
30'h0000016d: inst = 32'h13054512;
30'h0000016e: inst = 32'h23201500;
30'h0000016f: inst = 32'hb7801300;
30'h00000170: inst = 32'h93803039;
30'h00000171: inst = 32'h3705ff3f;
30'h00000172: inst = 32'h13058512;
30'h00000173: inst = 32'h23201500;
30'h00000174: inst = 32'hb7101000;
30'h00000175: inst = 32'h938030a1;
30'h00000176: inst = 32'h3705ff3f;
30'h00000177: inst = 32'h1305c512;
30'h00000178: inst = 32'h23201500;
30'h00000179: inst = 32'hb7102000;
30'h0000017a: inst = 32'h938030a9;
30'h0000017b: inst = 32'h3705ff3f;
30'h0000017c: inst = 32'h13050513;
30'h0000017d: inst = 32'h23201500;
30'h0000017e: inst = 32'h930070bb;
30'h0000017f: inst = 32'h3705ff3f;
30'h00000180: inst = 32'h13054513;
30'h00000181: inst = 32'h23201500;
30'h00000182: inst = 32'hb7505a59;
30'h00000183: inst = 32'h93803066;
30'h00000184: inst = 32'h3705ff3f;
30'h00000185: inst = 32'h13058513;
30'h00000186: inst = 32'h23201500;
30'h00000187: inst = 32'hb7d05b59;
30'h00000188: inst = 32'h93803046;
30'h00000189: inst = 32'h3705ff3f;
30'h0000018a: inst = 32'h1305c513;
30'h0000018b: inst = 32'h23201500;
30'h0000018c: inst = 32'hb7507a01;
30'h0000018d: inst = 32'h93803046;
30'h0000018e: inst = 32'h3705ff3f;
30'h0000018f: inst = 32'h13050514;
30'h00000190: inst = 32'h23201500;
30'h00000191: inst = 32'hb700c04d;
30'h00000192: inst = 32'h9380f006;
30'h00000193: inst = 32'h3705ff3f;
30'h00000194: inst = 32'h13054514;
30'h00000195: inst = 32'h23201500;
30'h00000196: inst = 32'hb7102006;
30'h00000197: inst = 32'h938030f9;
30'h00000198: inst = 32'h3705ff3f;
30'h00000199: inst = 32'h13058514;
30'h0000019a: inst = 32'h23201500;
30'h0000019b: inst = 32'hb7801300;
30'h0000019c: inst = 32'h93803039;
30'h0000019d: inst = 32'h3705ff3f;
30'h0000019e: inst = 32'h1305c514;
30'h0000019f: inst = 32'h23201500;
30'h000001a0: inst = 32'hb7101000;
30'h000001a1: inst = 32'h938030a1;
30'h000001a2: inst = 32'h3705ff3f;
30'h000001a3: inst = 32'h13050515;
30'h000001a4: inst = 32'h23201500;
30'h000001a5: inst = 32'hb7102000;
30'h000001a6: inst = 32'h938030a9;
30'h000001a7: inst = 32'h3705ff3f;
30'h000001a8: inst = 32'h13054515;
30'h000001a9: inst = 32'h23201500;
30'h000001aa: inst = 32'h930070bb;
30'h000001ab: inst = 32'h3705ff3f;
30'h000001ac: inst = 32'h13058515;
30'h000001ad: inst = 32'h23201500;
30'h000001ae: inst = 32'hb7707a57;
30'h000001af: inst = 32'h93803046;
30'h000001b0: inst = 32'h3705ff3f;
30'h000001b1: inst = 32'h1305c515;
30'h000001b2: inst = 32'h23201500;
30'h000001b3: inst = 32'hb7705a57;
30'h000001b4: inst = 32'h93803026;
30'h000001b5: inst = 32'h3705ff3f;
30'h000001b6: inst = 32'h13050516;
30'h000001b7: inst = 32'h23201500;
30'h000001b8: inst = 32'hb7705057;
30'h000001b9: inst = 32'h93803006;
30'h000001ba: inst = 32'h3705ff3f;
30'h000001bb: inst = 32'h13054516;
30'h000001bc: inst = 32'h23201500;
30'h000001bd: inst = 32'hb7f05b01;
30'h000001be: inst = 32'h93803046;
30'h000001bf: inst = 32'h3705ff3f;
30'h000001c0: inst = 32'h13058516;
30'h000001c1: inst = 32'h23201500;
30'h000001c2: inst = 32'hb700404b;
30'h000001c3: inst = 32'h9380f006;
30'h000001c4: inst = 32'h3705ff3f;
30'h000001c5: inst = 32'h1305c516;
30'h000001c6: inst = 32'h23201500;
30'h000001c7: inst = 32'hb7103006;
30'h000001c8: inst = 32'h938030f9;
30'h000001c9: inst = 32'h3705ff3f;
30'h000001ca: inst = 32'h13050517;
30'h000001cb: inst = 32'h23201500;
30'h000001cc: inst = 32'hb7801300;
30'h000001cd: inst = 32'h93803039;
30'h000001ce: inst = 32'h3705ff3f;
30'h000001cf: inst = 32'h13054517;
30'h000001d0: inst = 32'h23201500;
30'h000001d1: inst = 32'hb710f00f;
30'h000001d2: inst = 32'h938030a1;
30'h000001d3: inst = 32'h3705ff3f;
30'h000001d4: inst = 32'h13058517;
30'h000001d5: inst = 32'h23201500;
30'h000001d6: inst = 32'hb7204a01;
30'h000001d7: inst = 32'h938030a9;
30'h000001d8: inst = 32'h3705ff3f;
30'h000001d9: inst = 32'h1305c517;
30'h000001da: inst = 32'h23201500;
30'h000001db: inst = 32'hb710f00f;
30'h000001dc: inst = 32'h938070bb;
30'h000001dd: inst = 32'h3705ff3f;
30'h000001de: inst = 32'h13050518;
30'h000001df: inst = 32'h23201500;
30'h000001e0: inst = 32'hb7a05b49;
30'h000001e1: inst = 32'h938030e6;
30'h000001e2: inst = 32'h3705ff3f;
30'h000001e3: inst = 32'h13054518;
30'h000001e4: inst = 32'h23201500;
30'h000001e5: inst = 32'hb7104006;
30'h000001e6: inst = 32'h938030f9;
30'h000001e7: inst = 32'h3705ff3f;
30'h000001e8: inst = 32'h13058518;
30'h000001e9: inst = 32'h23201500;
30'h000001ea: inst = 32'hb7801300;
30'h000001eb: inst = 32'h93803039;
30'h000001ec: inst = 32'h3705ff3f;
30'h000001ed: inst = 32'h1305c518;
30'h000001ee: inst = 32'h23201500;
30'h000001ef: inst = 32'h930070c3;
30'h000001f0: inst = 32'h3705ff3f;
30'h000001f1: inst = 32'h13050519;
30'h000001f2: inst = 32'h23201500;
30'h000001f3: inst = 32'hb770fcff;
30'h000001f4: inst = 32'h938030c1;
30'h000001f5: inst = 32'h3705ff3f;
30'h000001f6: inst = 32'h13054519;
30'h000001f7: inst = 32'h23201500;
30'h000001f8: inst = 32'hb7100080;
30'h000001f9: inst = 32'h938070bb;
30'h000001fa: inst = 32'h3705ff3f;
30'h000001fb: inst = 32'h13058519;
30'h000001fc: inst = 32'h23201500;
30'h000001fd: inst = 32'hb7e0fb41;
30'h000001fe: inst = 32'h938030b9;
30'h000001ff: inst = 32'h3705ff3f;
30'h00000200: inst = 32'h1305c519;
30'h00000201: inst = 32'h23201500;
30'h00000202: inst = 32'hb7107c49;
30'h00000203: inst = 32'h93803006;
30'h00000204: inst = 32'h3705ff3f;
30'h00000205: inst = 32'h1305051a;
30'h00000206: inst = 32'h23201500;
30'h00000207: inst = 32'hb7105006;
30'h00000208: inst = 32'h938030f9;
30'h00000209: inst = 32'h3705ff3f;
30'h0000020a: inst = 32'h1305451a;
30'h0000020b: inst = 32'h23201500;
30'h0000020c: inst = 32'hb7801300;
30'h0000020d: inst = 32'h93803039;
30'h0000020e: inst = 32'h3705ff3f;
30'h0000020f: inst = 32'h1305851a;
30'h00000210: inst = 32'h23201500;
30'h00000211: inst = 32'hb7000010;
30'h00000212: inst = 32'h93807053;
30'h00000213: inst = 32'h3705ff3f;
30'h00000214: inst = 32'h1305c51a;
30'h00000215: inst = 32'h23201500;
30'h00000216: inst = 32'hb7506587;
30'h00000217: inst = 32'h938070ab;
30'h00000218: inst = 32'h3705ff3f;
30'h00000219: inst = 32'h1305051b;
30'h0000021a: inst = 32'h23201500;
30'h0000021b: inst = 32'hb7f01a32;
30'h0000021c: inst = 32'h938030a9;
30'h0000021d: inst = 32'h3705ff3f;
30'h0000021e: inst = 32'h1305451b;
30'h0000021f: inst = 32'h23201500;
30'h00000220: inst = 32'hb7205501;
30'h00000221: inst = 32'h93803002;
30'h00000222: inst = 32'h3705ff3f;
30'h00000223: inst = 32'h1305851b;
30'h00000224: inst = 32'h23201500;
30'h00000225: inst = 32'hb7100500;
30'h00000226: inst = 32'h938030b0;
30'h00000227: inst = 32'h3705ff3f;
30'h00000228: inst = 32'h1305c51b;
30'h00000229: inst = 32'h23201500;
30'h0000022a: inst = 32'hb7101002;
30'h0000022b: inst = 32'h938030c1;
30'h0000022c: inst = 32'h3705ff3f;
30'h0000022d: inst = 32'h1305051c;
30'h0000022e: inst = 32'h23201500;
30'h0000022f: inst = 32'hb7208b45;
30'h00000230: inst = 32'h938030e6;
30'h00000231: inst = 32'h3705ff3f;
30'h00000232: inst = 32'h1305451c;
30'h00000233: inst = 32'h23201500;
30'h00000234: inst = 32'hb7101500;
30'h00000235: inst = 32'h938030b0;
30'h00000236: inst = 32'h3705ff3f;
30'h00000237: inst = 32'h1305851c;
30'h00000238: inst = 32'h23201500;
30'h00000239: inst = 32'hb7103004;
30'h0000023a: inst = 32'h938030c1;
30'h0000023b: inst = 32'h3705ff3f;
30'h0000023c: inst = 32'h1305c51c;
30'h0000023d: inst = 32'h23201500;
30'h0000023e: inst = 32'hb7208b45;
30'h0000023f: inst = 32'h93803086;
30'h00000240: inst = 32'h3705ff3f;
30'h00000241: inst = 32'h1305051d;
30'h00000242: inst = 32'h23201500;
30'h00000243: inst = 32'hb7102500;
30'h00000244: inst = 32'h938030b0;
30'h00000245: inst = 32'h3705ff3f;
30'h00000246: inst = 32'h1305451d;
30'h00000247: inst = 32'h23201500;
30'h00000248: inst = 32'hb7105006;
30'h00000249: inst = 32'h938030c1;
30'h0000024a: inst = 32'h3705ff3f;
30'h0000024b: inst = 32'h1305851d;
30'h0000024c: inst = 32'h23201500;
30'h0000024d: inst = 32'hb7108b45;
30'h0000024e: inst = 32'h93803026;
30'h0000024f: inst = 32'h3705ff3f;
30'h00000250: inst = 32'h1305c51d;
30'h00000251: inst = 32'h23201500;
30'h00000252: inst = 32'hb7103500;
30'h00000253: inst = 32'h938030b0;
30'h00000254: inst = 32'h3705ff3f;
30'h00000255: inst = 32'h1305051e;
30'h00000256: inst = 32'h23201500;
30'h00000257: inst = 32'hb7100087;
30'h00000258: inst = 32'h938070c3;
30'h00000259: inst = 32'h3705ff3f;
30'h0000025a: inst = 32'h1305451e;
30'h0000025b: inst = 32'h23201500;
30'h0000025c: inst = 32'hb7608c41;
30'h0000025d: inst = 32'h938030c1;
30'h0000025e: inst = 32'h3705ff3f;
30'h0000025f: inst = 32'h1305851e;
30'h00000260: inst = 32'h23201500;
30'h00000261: inst = 32'hb7208b43;
30'h00000262: inst = 32'h938030a6;
30'h00000263: inst = 32'h3705ff3f;
30'h00000264: inst = 32'h1305c51e;
30'h00000265: inst = 32'h23201500;
30'h00000266: inst = 32'hb7106006;
30'h00000267: inst = 32'h938030f9;
30'h00000268: inst = 32'h3705ff3f;
30'h00000269: inst = 32'h1305051f;
30'h0000026a: inst = 32'h23201500;
30'h0000026b: inst = 32'hb7801300;
30'h0000026c: inst = 32'h93803039;
30'h0000026d: inst = 32'h3705ff3f;
30'h0000026e: inst = 32'h1305451f;
30'h0000026f: inst = 32'h23201500;
30'h00000270: inst = 32'hb7000010;
30'h00000271: inst = 32'h93807053;
30'h00000272: inst = 32'h3705ff3f;
30'h00000273: inst = 32'h1305851f;
30'h00000274: inst = 32'h23201500;
30'h00000275: inst = 32'hb710efcd;
30'h00000276: inst = 32'h938070d3;
30'h00000277: inst = 32'h3705ff3f;
30'h00000278: inst = 32'h1305c51f;
30'h00000279: inst = 32'h23201500;
30'h0000027a: inst = 32'hb7600d01;
30'h0000027b: inst = 32'h938030d1;
30'h0000027c: inst = 32'h3705ff3f;
30'h0000027d: inst = 32'h13050520;
30'h0000027e: inst = 32'h23201500;
30'h0000027f: inst = 32'hb710ab89;
30'h00000280: inst = 32'h938070a3;
30'h00000281: inst = 32'h3705ff3f;
30'h00000282: inst = 32'h13054520;
30'h00000283: inst = 32'h23201500;
30'h00000284: inst = 32'hb7104d01;
30'h00000285: inst = 32'h9380309b;
30'h00000286: inst = 32'h3705ff3f;
30'h00000287: inst = 32'h13058520;
30'h00000288: inst = 32'h23201500;
30'h00000289: inst = 32'hb7203501;
30'h0000028a: inst = 32'h93803002;
30'h0000028b: inst = 32'h3705ff3f;
30'h0000028c: inst = 32'h1305c520;
30'h0000028d: inst = 32'h23201500;
30'h0000028e: inst = 32'hb7200500;
30'h0000028f: inst = 32'h93803078;
30'h00000290: inst = 32'h3705ff3f;
30'h00000291: inst = 32'h13050521;
30'h00000292: inst = 32'h23201500;
30'h00000293: inst = 32'hb7100500;
30'h00000294: inst = 32'h938030b0;
30'h00000295: inst = 32'h3705ff3f;
30'h00000296: inst = 32'h13054521;
30'h00000297: inst = 32'h23201500;
30'h00000298: inst = 32'hb71000ef;
30'h00000299: inst = 32'h938070c3;
30'h0000029a: inst = 32'h3705ff3f;
30'h0000029b: inst = 32'h13058521;
30'h0000029c: inst = 32'h23201500;
30'h0000029d: inst = 32'hb7608c41;
30'h0000029e: inst = 32'h938030c1;
30'h0000029f: inst = 32'h3705ff3f;
30'h000002a0: inst = 32'h1305c521;
30'h000002a1: inst = 32'h23201500;
30'h000002a2: inst = 32'hb7108b41;
30'h000002a3: inst = 32'h93803006;
30'h000002a4: inst = 32'h3705ff3f;
30'h000002a5: inst = 32'h13050522;
30'h000002a6: inst = 32'h23201500;
30'h000002a7: inst = 32'hb7101500;
30'h000002a8: inst = 32'h938030b0;
30'h000002a9: inst = 32'h3705ff3f;
30'h000002aa: inst = 32'h13054522;
30'h000002ab: inst = 32'h23201500;
30'h000002ac: inst = 32'hb71000cd;
30'h000002ad: inst = 32'h938070c3;
30'h000002ae: inst = 32'h3705ff3f;
30'h000002af: inst = 32'h13058522;
30'h000002b0: inst = 32'h23201500;
30'h000002b1: inst = 32'hb7608c41;
30'h000002b2: inst = 32'h938030c1;
30'h000002b3: inst = 32'h3705ff3f;
30'h000002b4: inst = 32'h1305c522;
30'h000002b5: inst = 32'h23201500;
30'h000002b6: inst = 32'hb7208b3f;
30'h000002b7: inst = 32'h93803086;
30'h000002b8: inst = 32'h3705ff3f;
30'h000002b9: inst = 32'h13050523;
30'h000002ba: inst = 32'h23201500;
30'h000002bb: inst = 32'hb7102500;
30'h000002bc: inst = 32'h938030b0;
30'h000002bd: inst = 32'h3705ff3f;
30'h000002be: inst = 32'h13054523;
30'h000002bf: inst = 32'h23201500;
30'h000002c0: inst = 32'hb71000ab;
30'h000002c1: inst = 32'h938070c3;
30'h000002c2: inst = 32'h3705ff3f;
30'h000002c3: inst = 32'h13058523;
30'h000002c4: inst = 32'h23201500;
30'h000002c5: inst = 32'hb7608c41;
30'h000002c6: inst = 32'h938030c1;
30'h000002c7: inst = 32'h3705ff3f;
30'h000002c8: inst = 32'h1305c523;
30'h000002c9: inst = 32'h23201500;
30'h000002ca: inst = 32'hb7108b3f;
30'h000002cb: inst = 32'h93803006;
30'h000002cc: inst = 32'h3705ff3f;
30'h000002cd: inst = 32'h13050524;
30'h000002ce: inst = 32'h23201500;
30'h000002cf: inst = 32'hb7300500;
30'h000002d0: inst = 32'h938030c8;
30'h000002d1: inst = 32'h3705ff3f;
30'h000002d2: inst = 32'h13054524;
30'h000002d3: inst = 32'h23201500;
30'h000002d4: inst = 32'hb7103500;
30'h000002d5: inst = 32'h938030b0;
30'h000002d6: inst = 32'h3705ff3f;
30'h000002d7: inst = 32'h13058524;
30'h000002d8: inst = 32'h23201500;
30'h000002d9: inst = 32'hb7100089;
30'h000002da: inst = 32'h938070c3;
30'h000002db: inst = 32'h3705ff3f;
30'h000002dc: inst = 32'h1305c524;
30'h000002dd: inst = 32'h23201500;
30'h000002de: inst = 32'hb7608c41;
30'h000002df: inst = 32'h938030c1;
30'h000002e0: inst = 32'h3705ff3f;
30'h000002e1: inst = 32'h13050525;
30'h000002e2: inst = 32'h23201500;
30'h000002e3: inst = 32'hb7108b3d;
30'h000002e4: inst = 32'h93803066;
30'h000002e5: inst = 32'h3705ff3f;
30'h000002e6: inst = 32'h13054525;
30'h000002e7: inst = 32'h23201500;
30'h000002e8: inst = 32'hb7107006;
30'h000002e9: inst = 32'h938030f9;
30'h000002ea: inst = 32'h3705ff3f;
30'h000002eb: inst = 32'h13058525;
30'h000002ec: inst = 32'h23201500;
30'h000002ed: inst = 32'hb7801300;
30'h000002ee: inst = 32'h93803039;
30'h000002ef: inst = 32'h3705ff3f;
30'h000002f0: inst = 32'h1305c525;
30'h000002f1: inst = 32'h23201500;
30'h000002f2: inst = 32'hb7000010;
30'h000002f3: inst = 32'h93807053;
30'h000002f4: inst = 32'h3705ff3f;
30'h000002f5: inst = 32'h13050526;
30'h000002f6: inst = 32'h23201500;
30'h000002f7: inst = 32'hb710efcd;
30'h000002f8: inst = 32'h938070d3;
30'h000002f9: inst = 32'h3705ff3f;
30'h000002fa: inst = 32'h13054526;
30'h000002fb: inst = 32'h23201500;
30'h000002fc: inst = 32'hb7600d01;
30'h000002fd: inst = 32'h938030d1;
30'h000002fe: inst = 32'h3705ff3f;
30'h000002ff: inst = 32'h13058526;
30'h00000300: inst = 32'h23201500;
30'h00000301: inst = 32'hb710ab89;
30'h00000302: inst = 32'h938070a3;
30'h00000303: inst = 32'h3705ff3f;
30'h00000304: inst = 32'h1305c526;
30'h00000305: inst = 32'h23201500;
30'h00000306: inst = 32'hb7104d01;
30'h00000307: inst = 32'h9380309b;
30'h00000308: inst = 32'h3705ff3f;
30'h00000309: inst = 32'h13050527;
30'h0000030a: inst = 32'h23201500;
30'h0000030b: inst = 32'hb7203501;
30'h0000030c: inst = 32'h93803002;
30'h0000030d: inst = 32'h3705ff3f;
30'h0000030e: inst = 32'h13054527;
30'h0000030f: inst = 32'h23201500;
30'h00000310: inst = 32'hb7200500;
30'h00000311: inst = 32'h93803078;
30'h00000312: inst = 32'h3705ff3f;
30'h00000313: inst = 32'h13058527;
30'h00000314: inst = 32'h23201500;
30'h00000315: inst = 32'hb7200500;
30'h00000316: inst = 32'h938030b0;
30'h00000317: inst = 32'h3705ff3f;
30'h00000318: inst = 32'h1305c527;
30'h00000319: inst = 32'h23201500;
30'h0000031a: inst = 32'hb710efcd;
30'h0000031b: inst = 32'h938070c3;
30'h0000031c: inst = 32'h3705ff3f;
30'h0000031d: inst = 32'h13050528;
30'h0000031e: inst = 32'h23201500;
30'h0000031f: inst = 32'hb7600c41;
30'h00000320: inst = 32'h938030c1;
30'h00000321: inst = 32'h3705ff3f;
30'h00000322: inst = 32'h13054528;
30'h00000323: inst = 32'h23201500;
30'h00000324: inst = 32'hb7208b39;
30'h00000325: inst = 32'h938030c6;
30'h00000326: inst = 32'h3705ff3f;
30'h00000327: inst = 32'h13058528;
30'h00000328: inst = 32'h23201500;
30'h00000329: inst = 32'hb7202500;
30'h0000032a: inst = 32'h938030b0;
30'h0000032b: inst = 32'h3705ff3f;
30'h0000032c: inst = 32'h1305c528;
30'h0000032d: inst = 32'h23201500;
30'h0000032e: inst = 32'hb710ab89;
30'h0000032f: inst = 32'h938070c3;
30'h00000330: inst = 32'h3705ff3f;
30'h00000331: inst = 32'h13050529;
30'h00000332: inst = 32'h23201500;
30'h00000333: inst = 32'hb7600c41;
30'h00000334: inst = 32'h938030c1;
30'h00000335: inst = 32'h3705ff3f;
30'h00000336: inst = 32'h13054529;
30'h00000337: inst = 32'h23201500;
30'h00000338: inst = 32'hb7108b39;
30'h00000339: inst = 32'h93803046;
30'h0000033a: inst = 32'h3705ff3f;
30'h0000033b: inst = 32'h13058529;
30'h0000033c: inst = 32'h23201500;
30'h0000033d: inst = 32'hb7108006;
30'h0000033e: inst = 32'h938030f9;
30'h0000033f: inst = 32'h3705ff3f;
30'h00000340: inst = 32'h1305c529;
30'h00000341: inst = 32'h23201500;
30'h00000342: inst = 32'hb7801300;
30'h00000343: inst = 32'h93803039;
30'h00000344: inst = 32'h3705ff3f;
30'h00000345: inst = 32'h1305052a;
30'h00000346: inst = 32'h23201500;
30'h00000347: inst = 32'hb7000010;
30'h00000348: inst = 32'h93807053;
30'h00000349: inst = 32'h3705ff3f;
30'h0000034a: inst = 32'h1305452a;
30'h0000034b: inst = 32'h23201500;
30'h0000034c: inst = 32'hb7102143;
30'h0000034d: inst = 32'h938070d3;
30'h0000034e: inst = 32'h3705ff3f;
30'h0000034f: inst = 32'h1305852a;
30'h00000350: inst = 32'h23201500;
30'h00000351: inst = 32'hb7600d01;
30'h00000352: inst = 32'h938030d1;
30'h00000353: inst = 32'h3705ff3f;
30'h00000354: inst = 32'h1305c52a;
30'h00000355: inst = 32'h23201500;
30'h00000356: inst = 32'hb7106587;
30'h00000357: inst = 32'h938070a3;
30'h00000358: inst = 32'h3705ff3f;
30'h00000359: inst = 32'h1305052b;
30'h0000035a: inst = 32'h23201500;
30'h0000035b: inst = 32'hb7104d01;
30'h0000035c: inst = 32'h9380309b;
30'h0000035d: inst = 32'h3705ff3f;
30'h0000035e: inst = 32'h1305452b;
30'h0000035f: inst = 32'h23201500;
30'h00000360: inst = 32'hb7203501;
30'h00000361: inst = 32'h93803002;
30'h00000362: inst = 32'h3705ff3f;
30'h00000363: inst = 32'h1305852b;
30'h00000364: inst = 32'h23201500;
30'h00000365: inst = 32'hb7200500;
30'h00000366: inst = 32'h93803078;
30'h00000367: inst = 32'h3705ff3f;
30'h00000368: inst = 32'h1305c52b;
30'h00000369: inst = 32'h23201500;
30'h0000036a: inst = 32'hb7200500;
30'h0000036b: inst = 32'h938030b0;
30'h0000036c: inst = 32'h3705ff3f;
30'h0000036d: inst = 32'h1305052c;
30'h0000036e: inst = 32'h23201500;
30'h0000036f: inst = 32'hb7102143;
30'h00000370: inst = 32'h938070c3;
30'h00000371: inst = 32'h3705ff3f;
30'h00000372: inst = 32'h1305452c;
30'h00000373: inst = 32'h23201500;
30'h00000374: inst = 32'hb7600c41;
30'h00000375: inst = 32'h938030c1;
30'h00000376: inst = 32'h3705ff3f;
30'h00000377: inst = 32'h1305852c;
30'h00000378: inst = 32'h23201500;
30'h00000379: inst = 32'hb7208b35;
30'h0000037a: inst = 32'h938030a6;
30'h0000037b: inst = 32'h3705ff3f;
30'h0000037c: inst = 32'h1305c52c;
30'h0000037d: inst = 32'h23201500;
30'h0000037e: inst = 32'hb7202500;
30'h0000037f: inst = 32'h938030b0;
30'h00000380: inst = 32'h3705ff3f;
30'h00000381: inst = 32'h1305052d;
30'h00000382: inst = 32'h23201500;
30'h00000383: inst = 32'hb7106587;
30'h00000384: inst = 32'h938070c3;
30'h00000385: inst = 32'h3705ff3f;
30'h00000386: inst = 32'h1305452d;
30'h00000387: inst = 32'h23201500;
30'h00000388: inst = 32'hb7600c41;
30'h00000389: inst = 32'h938030c1;
30'h0000038a: inst = 32'h3705ff3f;
30'h0000038b: inst = 32'h1305852d;
30'h0000038c: inst = 32'h23201500;
30'h0000038d: inst = 32'hb7108b35;
30'h0000038e: inst = 32'h93803026;
30'h0000038f: inst = 32'h3705ff3f;
30'h00000390: inst = 32'h1305c52d;
30'h00000391: inst = 32'h23201500;
30'h00000392: inst = 32'hb7109006;
30'h00000393: inst = 32'h938030f9;
30'h00000394: inst = 32'h3705ff3f;
30'h00000395: inst = 32'h1305052e;
30'h00000396: inst = 32'h23201500;
30'h00000397: inst = 32'hb7801300;
30'h00000398: inst = 32'h93803039;
30'h00000399: inst = 32'h3705ff3f;
30'h0000039a: inst = 32'h1305452e;
30'h0000039b: inst = 32'h23201500;
30'h0000039c: inst = 32'hb7000010;
30'h0000039d: inst = 32'h93807053;
30'h0000039e: inst = 32'h3705ff3f;
30'h0000039f: inst = 32'h1305852e;
30'h000003a0: inst = 32'h23201500;
30'h000003a1: inst = 32'hb7102143;
30'h000003a2: inst = 32'h938070d3;
30'h000003a3: inst = 32'h3705ff3f;
30'h000003a4: inst = 32'h1305c52e;
30'h000003a5: inst = 32'h23201500;
30'h000003a6: inst = 32'hb7600d01;
30'h000003a7: inst = 32'h938030d1;
30'h000003a8: inst = 32'h3705ff3f;
30'h000003a9: inst = 32'h1305052f;
30'h000003aa: inst = 32'h23201500;
30'h000003ab: inst = 32'hb7106587;
30'h000003ac: inst = 32'h938070a3;
30'h000003ad: inst = 32'h3705ff3f;
30'h000003ae: inst = 32'h1305452f;
30'h000003af: inst = 32'h23201500;
30'h000003b0: inst = 32'hb7104d01;
30'h000003b1: inst = 32'h9380309b;
30'h000003b2: inst = 32'h3705ff3f;
30'h000003b3: inst = 32'h1305852f;
30'h000003b4: inst = 32'h23201500;
30'h000003b5: inst = 32'hb7203501;
30'h000003b6: inst = 32'h93803002;
30'h000003b7: inst = 32'h3705ff3f;
30'h000003b8: inst = 32'h1305c52f;
30'h000003b9: inst = 32'h23201500;
30'h000003ba: inst = 32'hb7200500;
30'h000003bb: inst = 32'h93803078;
30'h000003bc: inst = 32'h3705ff3f;
30'h000003bd: inst = 32'h13050530;
30'h000003be: inst = 32'h23201500;
30'h000003bf: inst = 32'hb7a03731;
30'h000003c0: inst = 32'h938030e6;
30'h000003c1: inst = 32'h3705ff3f;
30'h000003c2: inst = 32'h13054530;
30'h000003c3: inst = 32'h23201500;
30'h000003c4: inst = 32'hb710a006;
30'h000003c5: inst = 32'h938030f9;
30'h000003c6: inst = 32'h3705ff3f;
30'h000003c7: inst = 32'h13058530;
30'h000003c8: inst = 32'h23201500;
30'h000003c9: inst = 32'hb7801300;
30'h000003ca: inst = 32'h93803039;
30'h000003cb: inst = 32'h3705ff3f;
30'h000003cc: inst = 32'h1305c530;
30'h000003cd: inst = 32'h23201500;
30'h000003ce: inst = 32'hb7000010;
30'h000003cf: inst = 32'h93807053;
30'h000003d0: inst = 32'h3705ff3f;
30'h000003d1: inst = 32'h13050531;
30'h000003d2: inst = 32'h23201500;
30'h000003d3: inst = 32'hb7506587;
30'h000003d4: inst = 32'h938070ab;
30'h000003d5: inst = 32'h3705ff3f;
30'h000003d6: inst = 32'h13054531;
30'h000003d7: inst = 32'h23201500;
30'h000003d8: inst = 32'hb7f01a32;
30'h000003d9: inst = 32'h938030a9;
30'h000003da: inst = 32'h3705ff3f;
30'h000003db: inst = 32'h13058531;
30'h000003dc: inst = 32'h23201500;
30'h000003dd: inst = 32'hb7205501;
30'h000003de: inst = 32'h93803002;
30'h000003df: inst = 32'h3705ff3f;
30'h000003e0: inst = 32'h1305c531;
30'h000003e1: inst = 32'h23201500;
30'h000003e2: inst = 32'hb7500500;
30'h000003e3: inst = 32'h938030b0;
30'h000003e4: inst = 32'h3705ff3f;
30'h000003e5: inst = 32'h13050532;
30'h000003e6: inst = 32'h23201500;
30'h000003e7: inst = 32'hb7101002;
30'h000003e8: inst = 32'h938030c1;
30'h000003e9: inst = 32'h3705ff3f;
30'h000003ea: inst = 32'h13054532;
30'h000003eb: inst = 32'h23201500;
30'h000003ec: inst = 32'hb7208b2f;
30'h000003ed: inst = 32'h938030c6;
30'h000003ee: inst = 32'h3705ff3f;
30'h000003ef: inst = 32'h13058532;
30'h000003f0: inst = 32'h23201500;
30'h000003f1: inst = 32'hb7501500;
30'h000003f2: inst = 32'h938030b0;
30'h000003f3: inst = 32'h3705ff3f;
30'h000003f4: inst = 32'h1305c532;
30'h000003f5: inst = 32'h23201500;
30'h000003f6: inst = 32'hb7103004;
30'h000003f7: inst = 32'h938030c1;
30'h000003f8: inst = 32'h3705ff3f;
30'h000003f9: inst = 32'h13050533;
30'h000003fa: inst = 32'h23201500;
30'h000003fb: inst = 32'hb7108b2f;
30'h000003fc: inst = 32'h93803066;
30'h000003fd: inst = 32'h3705ff3f;
30'h000003fe: inst = 32'h13054533;
30'h000003ff: inst = 32'h23201500;
30'h00000400: inst = 32'hb7502500;
30'h00000401: inst = 32'h938030b0;
30'h00000402: inst = 32'h3705ff3f;
30'h00000403: inst = 32'h13058533;
30'h00000404: inst = 32'h23201500;
30'h00000405: inst = 32'hb7105006;
30'h00000406: inst = 32'h938030c1;
30'h00000407: inst = 32'h3705ff3f;
30'h00000408: inst = 32'h1305c533;
30'h00000409: inst = 32'h23201500;
30'h0000040a: inst = 32'hb7108b2f;
30'h0000040b: inst = 32'h93803006;
30'h0000040c: inst = 32'h3705ff3f;
30'h0000040d: inst = 32'h13050534;
30'h0000040e: inst = 32'h23201500;
30'h0000040f: inst = 32'hb7503500;
30'h00000410: inst = 32'h938030b0;
30'h00000411: inst = 32'h3705ff3f;
30'h00000412: inst = 32'h13054534;
30'h00000413: inst = 32'h23201500;
30'h00000414: inst = 32'hb7100087;
30'h00000415: inst = 32'h938070c3;
30'h00000416: inst = 32'h3705ff3f;
30'h00000417: inst = 32'h13058534;
30'h00000418: inst = 32'h23201500;
30'h00000419: inst = 32'hb7608c01;
30'h0000041a: inst = 32'h938030c1;
30'h0000041b: inst = 32'h3705ff3f;
30'h0000041c: inst = 32'h1305c534;
30'h0000041d: inst = 32'h23201500;
30'h0000041e: inst = 32'hb7208b2d;
30'h0000041f: inst = 32'h93803086;
30'h00000420: inst = 32'h3705ff3f;
30'h00000421: inst = 32'h13050535;
30'h00000422: inst = 32'h23201500;
30'h00000423: inst = 32'hb710b006;
30'h00000424: inst = 32'h938030f9;
30'h00000425: inst = 32'h3705ff3f;
30'h00000426: inst = 32'h13054535;
30'h00000427: inst = 32'h23201500;
30'h00000428: inst = 32'hb7801300;
30'h00000429: inst = 32'h93803039;
30'h0000042a: inst = 32'h3705ff3f;
30'h0000042b: inst = 32'h13058535;
30'h0000042c: inst = 32'h23201500;
30'h0000042d: inst = 32'hb7000010;
30'h0000042e: inst = 32'h93807053;
30'h0000042f: inst = 32'h3705ff3f;
30'h00000430: inst = 32'h1305c535;
30'h00000431: inst = 32'h23201500;
30'h00000432: inst = 32'hb710efcd;
30'h00000433: inst = 32'h938070d3;
30'h00000434: inst = 32'h3705ff3f;
30'h00000435: inst = 32'h13050536;
30'h00000436: inst = 32'h23201500;
30'h00000437: inst = 32'hb7600d01;
30'h00000438: inst = 32'h938030d1;
30'h00000439: inst = 32'h3705ff3f;
30'h0000043a: inst = 32'h13054536;
30'h0000043b: inst = 32'h23201500;
30'h0000043c: inst = 32'hb710ab89;
30'h0000043d: inst = 32'h938070a3;
30'h0000043e: inst = 32'h3705ff3f;
30'h0000043f: inst = 32'h13058536;
30'h00000440: inst = 32'h23201500;
30'h00000441: inst = 32'hb7104d01;
30'h00000442: inst = 32'h9380309b;
30'h00000443: inst = 32'h3705ff3f;
30'h00000444: inst = 32'h1305c536;
30'h00000445: inst = 32'h23201500;
30'h00000446: inst = 32'hb7203501;
30'h00000447: inst = 32'h93803002;
30'h00000448: inst = 32'h3705ff3f;
30'h00000449: inst = 32'h13050537;
30'h0000044a: inst = 32'h23201500;
30'h0000044b: inst = 32'hb7200500;
30'h0000044c: inst = 32'h93803078;
30'h0000044d: inst = 32'h3705ff3f;
30'h0000044e: inst = 32'h13054537;
30'h0000044f: inst = 32'h23201500;
30'h00000450: inst = 32'hb7500500;
30'h00000451: inst = 32'h938030b0;
30'h00000452: inst = 32'h3705ff3f;
30'h00000453: inst = 32'h13058537;
30'h00000454: inst = 32'h23201500;
30'h00000455: inst = 32'hb71000ef;
30'h00000456: inst = 32'h938070c3;
30'h00000457: inst = 32'h3705ff3f;
30'h00000458: inst = 32'h1305c537;
30'h00000459: inst = 32'h23201500;
30'h0000045a: inst = 32'hb7608c01;
30'h0000045b: inst = 32'h938030c1;
30'h0000045c: inst = 32'h3705ff3f;
30'h0000045d: inst = 32'h13050538;
30'h0000045e: inst = 32'h23201500;
30'h0000045f: inst = 32'hb7208b29;
30'h00000460: inst = 32'h938030e6;
30'h00000461: inst = 32'h3705ff3f;
30'h00000462: inst = 32'h13054538;
30'h00000463: inst = 32'h23201500;
30'h00000464: inst = 32'hb7501500;
30'h00000465: inst = 32'h938030b0;
30'h00000466: inst = 32'h3705ff3f;
30'h00000467: inst = 32'h13058538;
30'h00000468: inst = 32'h23201500;
30'h00000469: inst = 32'hb71000cd;
30'h0000046a: inst = 32'h938070c3;
30'h0000046b: inst = 32'h3705ff3f;
30'h0000046c: inst = 32'h1305c538;
30'h0000046d: inst = 32'h23201500;
30'h0000046e: inst = 32'hb7608c01;
30'h0000046f: inst = 32'h938030c1;
30'h00000470: inst = 32'h3705ff3f;
30'h00000471: inst = 32'h13050539;
30'h00000472: inst = 32'h23201500;
30'h00000473: inst = 32'hb7108b29;
30'h00000474: inst = 32'h93803066;
30'h00000475: inst = 32'h3705ff3f;
30'h00000476: inst = 32'h13054539;
30'h00000477: inst = 32'h23201500;
30'h00000478: inst = 32'hb7502500;
30'h00000479: inst = 32'h938030b0;
30'h0000047a: inst = 32'h3705ff3f;
30'h0000047b: inst = 32'h13058539;
30'h0000047c: inst = 32'h23201500;
30'h0000047d: inst = 32'hb71000ab;
30'h0000047e: inst = 32'h938070c3;
30'h0000047f: inst = 32'h3705ff3f;
30'h00000480: inst = 32'h1305c539;
30'h00000481: inst = 32'h23201500;
30'h00000482: inst = 32'hb7608c01;
30'h00000483: inst = 32'h938030c1;
30'h00000484: inst = 32'h3705ff3f;
30'h00000485: inst = 32'h1305053a;
30'h00000486: inst = 32'h23201500;
30'h00000487: inst = 32'hb7208b27;
30'h00000488: inst = 32'h938030e6;
30'h00000489: inst = 32'h3705ff3f;
30'h0000048a: inst = 32'h1305453a;
30'h0000048b: inst = 32'h23201500;
30'h0000048c: inst = 32'hb7503500;
30'h0000048d: inst = 32'h938030b0;
30'h0000048e: inst = 32'h3705ff3f;
30'h0000048f: inst = 32'h1305853a;
30'h00000490: inst = 32'h23201500;
30'h00000491: inst = 32'hb7100089;
30'h00000492: inst = 32'h938070c3;
30'h00000493: inst = 32'h3705ff3f;
30'h00000494: inst = 32'h1305c53a;
30'h00000495: inst = 32'h23201500;
30'h00000496: inst = 32'hb7608c01;
30'h00000497: inst = 32'h938030c1;
30'h00000498: inst = 32'h3705ff3f;
30'h00000499: inst = 32'h1305053b;
30'h0000049a: inst = 32'h23201500;
30'h0000049b: inst = 32'hb7108b27;
30'h0000049c: inst = 32'h93803066;
30'h0000049d: inst = 32'h3705ff3f;
30'h0000049e: inst = 32'h1305453b;
30'h0000049f: inst = 32'h23201500;
30'h000004a0: inst = 32'hb710c006;
30'h000004a1: inst = 32'h938030f9;
30'h000004a2: inst = 32'h3705ff3f;
30'h000004a3: inst = 32'h1305853b;
30'h000004a4: inst = 32'h23201500;
30'h000004a5: inst = 32'hb7801300;
30'h000004a6: inst = 32'h93803039;
30'h000004a7: inst = 32'h3705ff3f;
30'h000004a8: inst = 32'h1305c53b;
30'h000004a9: inst = 32'h23201500;
30'h000004aa: inst = 32'hb7000010;
30'h000004ab: inst = 32'h93807053;
30'h000004ac: inst = 32'h3705ff3f;
30'h000004ad: inst = 32'h1305053c;
30'h000004ae: inst = 32'h23201500;
30'h000004af: inst = 32'hb710efcd;
30'h000004b0: inst = 32'h938070d3;
30'h000004b1: inst = 32'h3705ff3f;
30'h000004b2: inst = 32'h1305453c;
30'h000004b3: inst = 32'h23201500;
30'h000004b4: inst = 32'hb7600d01;
30'h000004b5: inst = 32'h938030d1;
30'h000004b6: inst = 32'h3705ff3f;
30'h000004b7: inst = 32'h1305853c;
30'h000004b8: inst = 32'h23201500;
30'h000004b9: inst = 32'hb710ab89;
30'h000004ba: inst = 32'h938070a3;
30'h000004bb: inst = 32'h3705ff3f;
30'h000004bc: inst = 32'h1305c53c;
30'h000004bd: inst = 32'h23201500;
30'h000004be: inst = 32'hb7104d01;
30'h000004bf: inst = 32'h9380309b;
30'h000004c0: inst = 32'h3705ff3f;
30'h000004c1: inst = 32'h1305053d;
30'h000004c2: inst = 32'h23201500;
30'h000004c3: inst = 32'hb7203501;
30'h000004c4: inst = 32'h93803002;
30'h000004c5: inst = 32'h3705ff3f;
30'h000004c6: inst = 32'h1305453d;
30'h000004c7: inst = 32'h23201500;
30'h000004c8: inst = 32'hb7200500;
30'h000004c9: inst = 32'h93803078;
30'h000004ca: inst = 32'h3705ff3f;
30'h000004cb: inst = 32'h1305853d;
30'h000004cc: inst = 32'h23201500;
30'h000004cd: inst = 32'hb7600500;
30'h000004ce: inst = 32'h938030b0;
30'h000004cf: inst = 32'h3705ff3f;
30'h000004d0: inst = 32'h1305c53d;
30'h000004d1: inst = 32'h23201500;
30'h000004d2: inst = 32'hb710efcd;
30'h000004d3: inst = 32'h938070c3;
30'h000004d4: inst = 32'h3705ff3f;
30'h000004d5: inst = 32'h1305053e;
30'h000004d6: inst = 32'h23201500;
30'h000004d7: inst = 32'hb7600c01;
30'h000004d8: inst = 32'h938030c1;
30'h000004d9: inst = 32'h3705ff3f;
30'h000004da: inst = 32'h1305453e;
30'h000004db: inst = 32'h23201500;
30'h000004dc: inst = 32'hb7208b23;
30'h000004dd: inst = 32'h938030c6;
30'h000004de: inst = 32'h3705ff3f;
30'h000004df: inst = 32'h1305853e;
30'h000004e0: inst = 32'h23201500;
30'h000004e1: inst = 32'hb7602500;
30'h000004e2: inst = 32'h938030b0;
30'h000004e3: inst = 32'h3705ff3f;
30'h000004e4: inst = 32'h1305c53e;
30'h000004e5: inst = 32'h23201500;
30'h000004e6: inst = 32'hb710ab89;
30'h000004e7: inst = 32'h938070c3;
30'h000004e8: inst = 32'h3705ff3f;
30'h000004e9: inst = 32'h1305053f;
30'h000004ea: inst = 32'h23201500;
30'h000004eb: inst = 32'hb7600c01;
30'h000004ec: inst = 32'h938030c1;
30'h000004ed: inst = 32'h3705ff3f;
30'h000004ee: inst = 32'h1305453f;
30'h000004ef: inst = 32'h23201500;
30'h000004f0: inst = 32'hb7108b23;
30'h000004f1: inst = 32'h93803046;
30'h000004f2: inst = 32'h3705ff3f;
30'h000004f3: inst = 32'h1305853f;
30'h000004f4: inst = 32'h23201500;
30'h000004f5: inst = 32'hb710d006;
30'h000004f6: inst = 32'h938030f9;
30'h000004f7: inst = 32'h3705ff3f;
30'h000004f8: inst = 32'h1305c53f;
30'h000004f9: inst = 32'h23201500;
30'h000004fa: inst = 32'hb7801300;
30'h000004fb: inst = 32'h93803039;
30'h000004fc: inst = 32'h3705ff3f;
30'h000004fd: inst = 32'h13050540;
30'h000004fe: inst = 32'h23201500;
30'h000004ff: inst = 32'hb7000010;
30'h00000500: inst = 32'h93807053;
30'h00000501: inst = 32'h3705ff3f;
30'h00000502: inst = 32'h13054540;
30'h00000503: inst = 32'h23201500;
30'h00000504: inst = 32'hb7102143;
30'h00000505: inst = 32'h938070d3;
30'h00000506: inst = 32'h3705ff3f;
30'h00000507: inst = 32'h13058540;
30'h00000508: inst = 32'h23201500;
30'h00000509: inst = 32'hb7600d01;
30'h0000050a: inst = 32'h938030d1;
30'h0000050b: inst = 32'h3705ff3f;
30'h0000050c: inst = 32'h1305c540;
30'h0000050d: inst = 32'h23201500;
30'h0000050e: inst = 32'hb7106587;
30'h0000050f: inst = 32'h938070a3;
30'h00000510: inst = 32'h3705ff3f;
30'h00000511: inst = 32'h13050541;
30'h00000512: inst = 32'h23201500;
30'h00000513: inst = 32'hb7104d01;
30'h00000514: inst = 32'h9380309b;
30'h00000515: inst = 32'h3705ff3f;
30'h00000516: inst = 32'h13054541;
30'h00000517: inst = 32'h23201500;
30'h00000518: inst = 32'hb7203501;
30'h00000519: inst = 32'h93803002;
30'h0000051a: inst = 32'h3705ff3f;
30'h0000051b: inst = 32'h13058541;
30'h0000051c: inst = 32'h23201500;
30'h0000051d: inst = 32'hb7200500;
30'h0000051e: inst = 32'h93803078;
30'h0000051f: inst = 32'h3705ff3f;
30'h00000520: inst = 32'h1305c541;
30'h00000521: inst = 32'h23201500;
30'h00000522: inst = 32'hb7600500;
30'h00000523: inst = 32'h938030b0;
30'h00000524: inst = 32'h3705ff3f;
30'h00000525: inst = 32'h13050542;
30'h00000526: inst = 32'h23201500;
30'h00000527: inst = 32'hb7102143;
30'h00000528: inst = 32'h938070c3;
30'h00000529: inst = 32'h3705ff3f;
30'h0000052a: inst = 32'h13054542;
30'h0000052b: inst = 32'h23201500;
30'h0000052c: inst = 32'hb7600c01;
30'h0000052d: inst = 32'h938030c1;
30'h0000052e: inst = 32'h3705ff3f;
30'h0000052f: inst = 32'h13058542;
30'h00000530: inst = 32'h23201500;
30'h00000531: inst = 32'hb7208b1f;
30'h00000532: inst = 32'h938030a6;
30'h00000533: inst = 32'h3705ff3f;
30'h00000534: inst = 32'h1305c542;
30'h00000535: inst = 32'h23201500;
30'h00000536: inst = 32'hb7602500;
30'h00000537: inst = 32'h938030b0;
30'h00000538: inst = 32'h3705ff3f;
30'h00000539: inst = 32'h13050543;
30'h0000053a: inst = 32'h23201500;
30'h0000053b: inst = 32'hb7106587;
30'h0000053c: inst = 32'h938070c3;
30'h0000053d: inst = 32'h3705ff3f;
30'h0000053e: inst = 32'h13054543;
30'h0000053f: inst = 32'h23201500;
30'h00000540: inst = 32'hb7600c01;
30'h00000541: inst = 32'h938030c1;
30'h00000542: inst = 32'h3705ff3f;
30'h00000543: inst = 32'h13058543;
30'h00000544: inst = 32'h23201500;
30'h00000545: inst = 32'hb7108b1f;
30'h00000546: inst = 32'h93803026;
30'h00000547: inst = 32'h3705ff3f;
30'h00000548: inst = 32'h1305c543;
30'h00000549: inst = 32'h23201500;
30'h0000054a: inst = 32'hb710e006;
30'h0000054b: inst = 32'h938030f9;
30'h0000054c: inst = 32'h3705ff3f;
30'h0000054d: inst = 32'h13050544;
30'h0000054e: inst = 32'h23201500;
30'h0000054f: inst = 32'hb7801300;
30'h00000550: inst = 32'h93803039;
30'h00000551: inst = 32'h3705ff3f;
30'h00000552: inst = 32'h13054544;
30'h00000553: inst = 32'h23201500;
30'h00000554: inst = 32'hb7000010;
30'h00000555: inst = 32'h93807053;
30'h00000556: inst = 32'h3705ff3f;
30'h00000557: inst = 32'h13058544;
30'h00000558: inst = 32'h23201500;
30'h00000559: inst = 32'hb7102143;
30'h0000055a: inst = 32'h938070d3;
30'h0000055b: inst = 32'h3705ff3f;
30'h0000055c: inst = 32'h1305c544;
30'h0000055d: inst = 32'h23201500;
30'h0000055e: inst = 32'hb7600d01;
30'h0000055f: inst = 32'h938030d1;
30'h00000560: inst = 32'h3705ff3f;
30'h00000561: inst = 32'h13050545;
30'h00000562: inst = 32'h23201500;
30'h00000563: inst = 32'hb7106587;
30'h00000564: inst = 32'h938070a3;
30'h00000565: inst = 32'h3705ff3f;
30'h00000566: inst = 32'h13054545;
30'h00000567: inst = 32'h23201500;
30'h00000568: inst = 32'hb7104d01;
30'h00000569: inst = 32'h9380309b;
30'h0000056a: inst = 32'h3705ff3f;
30'h0000056b: inst = 32'h13058545;
30'h0000056c: inst = 32'h23201500;
30'h0000056d: inst = 32'hb7200500;
30'h0000056e: inst = 32'h93803002;
30'h0000056f: inst = 32'h3705ff3f;
30'h00000570: inst = 32'h1305c545;
30'h00000571: inst = 32'h23201500;
30'h00000572: inst = 32'hb7003501;
30'h00000573: inst = 32'h93803002;
30'h00000574: inst = 32'h3705ff3f;
30'h00000575: inst = 32'h13050546;
30'h00000576: inst = 32'h23201500;
30'h00000577: inst = 32'hb7100021;
30'h00000578: inst = 32'h938070c3;
30'h00000579: inst = 32'h3705ff3f;
30'h0000057a: inst = 32'h13054546;
30'h0000057b: inst = 32'h23201500;
30'h0000057c: inst = 32'hb7608c01;
30'h0000057d: inst = 32'h938030c1;
30'h0000057e: inst = 32'h3705ff3f;
30'h0000057f: inst = 32'h13058546;
30'h00000580: inst = 32'h23201500;
30'h00000581: inst = 32'hb7300500;
30'h00000582: inst = 32'h938030b0;
30'h00000583: inst = 32'h3705ff3f;
30'h00000584: inst = 32'h1305c546;
30'h00000585: inst = 32'h23201500;
30'h00000586: inst = 32'hb7208b1b;
30'h00000587: inst = 32'h93803086;
30'h00000588: inst = 32'h3705ff3f;
30'h00000589: inst = 32'h13050547;
30'h0000058a: inst = 32'h23201500;
30'h0000058b: inst = 32'hb7003501;
30'h0000058c: inst = 32'h9380300a;
30'h0000058d: inst = 32'h3705ff3f;
30'h0000058e: inst = 32'h13054547;
30'h0000058f: inst = 32'h23201500;
30'h00000590: inst = 32'hb7102121;
30'h00000591: inst = 32'h938070c3;
30'h00000592: inst = 32'h3705ff3f;
30'h00000593: inst = 32'h13058547;
30'h00000594: inst = 32'h23201500;
30'h00000595: inst = 32'hb7600c01;
30'h00000596: inst = 32'h938030c1;
30'h00000597: inst = 32'h3705ff3f;
30'h00000598: inst = 32'h1305c547;
30'h00000599: inst = 32'h23201500;
30'h0000059a: inst = 32'hb7300500;
30'h0000059b: inst = 32'h938030b0;
30'h0000059c: inst = 32'h3705ff3f;
30'h0000059d: inst = 32'h13050548;
30'h0000059e: inst = 32'h23201500;
30'h0000059f: inst = 32'hb7208b19;
30'h000005a0: inst = 32'h938030e6;
30'h000005a1: inst = 32'h3705ff3f;
30'h000005a2: inst = 32'h13054548;
30'h000005a3: inst = 32'h23201500;
30'h000005a4: inst = 32'hb7200500;
30'h000005a5: inst = 32'h93803002;
30'h000005a6: inst = 32'h3705ff3f;
30'h000005a7: inst = 32'h13058548;
30'h000005a8: inst = 32'h23201500;
30'h000005a9: inst = 32'hb7003501;
30'h000005aa: inst = 32'h93803012;
30'h000005ab: inst = 32'h3705ff3f;
30'h000005ac: inst = 32'h1305c548;
30'h000005ad: inst = 32'h23201500;
30'h000005ae: inst = 32'hb7102100;
30'h000005af: inst = 32'h938070c3;
30'h000005b0: inst = 32'h3705ff3f;
30'h000005b1: inst = 32'h13050549;
30'h000005b2: inst = 32'h23201500;
30'h000005b3: inst = 32'hb7300500;
30'h000005b4: inst = 32'h938030b0;
30'h000005b5: inst = 32'h3705ff3f;
30'h000005b6: inst = 32'h13054549;
30'h000005b7: inst = 32'h23201500;
30'h000005b8: inst = 32'hb7108b19;
30'h000005b9: inst = 32'h93803046;
30'h000005ba: inst = 32'h3705ff3f;
30'h000005bb: inst = 32'h13058549;
30'h000005bc: inst = 32'h23201500;
30'h000005bd: inst = 32'hb7003501;
30'h000005be: inst = 32'h9380301a;
30'h000005bf: inst = 32'h3705ff3f;
30'h000005c0: inst = 32'h1305c549;
30'h000005c1: inst = 32'h23201500;
30'h000005c2: inst = 32'hb7102121;
30'h000005c3: inst = 32'h938070c3;
30'h000005c4: inst = 32'h3705ff3f;
30'h000005c5: inst = 32'h1305054a;
30'h000005c6: inst = 32'h23201500;
30'h000005c7: inst = 32'hb7300500;
30'h000005c8: inst = 32'h938030b0;
30'h000005c9: inst = 32'h3705ff3f;
30'h000005ca: inst = 32'h1305454a;
30'h000005cb: inst = 32'h23201500;
30'h000005cc: inst = 32'hb7208b17;
30'h000005cd: inst = 32'h938030c6;
30'h000005ce: inst = 32'h3705ff3f;
30'h000005cf: inst = 32'h1305854a;
30'h000005d0: inst = 32'h23201500;
30'h000005d1: inst = 32'hb710e006;
30'h000005d2: inst = 32'h938030f9;
30'h000005d3: inst = 32'h3705ff3f;
30'h000005d4: inst = 32'h1305c54a;
30'h000005d5: inst = 32'h23201500;
30'h000005d6: inst = 32'hb7801300;
30'h000005d7: inst = 32'h93803039;
30'h000005d8: inst = 32'h3705ff3f;
30'h000005d9: inst = 32'h1305054b;
30'h000005da: inst = 32'h23201500;
30'h000005db: inst = 32'hb7000010;
30'h000005dc: inst = 32'h93807053;
30'h000005dd: inst = 32'h3705ff3f;
30'h000005de: inst = 32'h1305454b;
30'h000005df: inst = 32'h23201500;
30'h000005e0: inst = 32'hb7102143;
30'h000005e1: inst = 32'h938070d3;
30'h000005e2: inst = 32'h3705ff3f;
30'h000005e3: inst = 32'h1305854b;
30'h000005e4: inst = 32'h23201500;
30'h000005e5: inst = 32'hb7600d01;
30'h000005e6: inst = 32'h938030d1;
30'h000005e7: inst = 32'h3705ff3f;
30'h000005e8: inst = 32'h1305c54b;
30'h000005e9: inst = 32'h23201500;
30'h000005ea: inst = 32'hb7106587;
30'h000005eb: inst = 32'h938070a3;
30'h000005ec: inst = 32'h3705ff3f;
30'h000005ed: inst = 32'h1305054c;
30'h000005ee: inst = 32'h23201500;
30'h000005ef: inst = 32'hb7104d01;
30'h000005f0: inst = 32'h9380309b;
30'h000005f1: inst = 32'h3705ff3f;
30'h000005f2: inst = 32'h1305454c;
30'h000005f3: inst = 32'h23201500;
30'h000005f4: inst = 32'hb7200500;
30'h000005f5: inst = 32'h93803002;
30'h000005f6: inst = 32'h3705ff3f;
30'h000005f7: inst = 32'h1305854c;
30'h000005f8: inst = 32'h23201500;
30'h000005f9: inst = 32'hb7003501;
30'h000005fa: inst = 32'h93803002;
30'h000005fb: inst = 32'h3705ff3f;
30'h000005fc: inst = 32'h1305c54c;
30'h000005fd: inst = 32'h23201500;
30'h000005fe: inst = 32'hb7100021;
30'h000005ff: inst = 32'h938070c3;
30'h00000600: inst = 32'h3705ff3f;
30'h00000601: inst = 32'h1305054d;
30'h00000602: inst = 32'h23201500;
30'h00000603: inst = 32'hb7608c01;
30'h00000604: inst = 32'h938030c1;
30'h00000605: inst = 32'h3705ff3f;
30'h00000606: inst = 32'h1305454d;
30'h00000607: inst = 32'h23201500;
30'h00000608: inst = 32'hb7300500;
30'h00000609: inst = 32'h938030b0;
30'h0000060a: inst = 32'h3705ff3f;
30'h0000060b: inst = 32'h1305854d;
30'h0000060c: inst = 32'h23201500;
30'h0000060d: inst = 32'hb7108b15;
30'h0000060e: inst = 32'h93803026;
30'h0000060f: inst = 32'h3705ff3f;
30'h00000610: inst = 32'h1305c54d;
30'h00000611: inst = 32'h23201500;
30'h00000612: inst = 32'hb7003501;
30'h00000613: inst = 32'h9380300a;
30'h00000614: inst = 32'h3705ff3f;
30'h00000615: inst = 32'h1305054e;
30'h00000616: inst = 32'h23201500;
30'h00000617: inst = 32'hb7102121;
30'h00000618: inst = 32'h938070c3;
30'h00000619: inst = 32'h3705ff3f;
30'h0000061a: inst = 32'h1305454e;
30'h0000061b: inst = 32'h23201500;
30'h0000061c: inst = 32'hb7600c01;
30'h0000061d: inst = 32'h938030c1;
30'h0000061e: inst = 32'h3705ff3f;
30'h0000061f: inst = 32'h1305854e;
30'h00000620: inst = 32'h23201500;
30'h00000621: inst = 32'hb7300500;
30'h00000622: inst = 32'h938030b0;
30'h00000623: inst = 32'h3705ff3f;
30'h00000624: inst = 32'h1305c54e;
30'h00000625: inst = 32'h23201500;
30'h00000626: inst = 32'hb7208b13;
30'h00000627: inst = 32'h93803086;
30'h00000628: inst = 32'h3705ff3f;
30'h00000629: inst = 32'h1305054f;
30'h0000062a: inst = 32'h23201500;
30'h0000062b: inst = 32'hb7200500;
30'h0000062c: inst = 32'h93803002;
30'h0000062d: inst = 32'h3705ff3f;
30'h0000062e: inst = 32'h1305454f;
30'h0000062f: inst = 32'h23201500;
30'h00000630: inst = 32'hb7003501;
30'h00000631: inst = 32'h93803012;
30'h00000632: inst = 32'h3705ff3f;
30'h00000633: inst = 32'h1305854f;
30'h00000634: inst = 32'h23201500;
30'h00000635: inst = 32'hb7102100;
30'h00000636: inst = 32'h938070c3;
30'h00000637: inst = 32'h3705ff3f;
30'h00000638: inst = 32'h1305c54f;
30'h00000639: inst = 32'h23201500;
30'h0000063a: inst = 32'hb7300500;
30'h0000063b: inst = 32'h938030b0;
30'h0000063c: inst = 32'h3705ff3f;
30'h0000063d: inst = 32'h13050550;
30'h0000063e: inst = 32'h23201500;
30'h0000063f: inst = 32'hb7208b11;
30'h00000640: inst = 32'h938030e6;
30'h00000641: inst = 32'h3705ff3f;
30'h00000642: inst = 32'h13054550;
30'h00000643: inst = 32'h23201500;
30'h00000644: inst = 32'hb7003501;
30'h00000645: inst = 32'h9380301a;
30'h00000646: inst = 32'h3705ff3f;
30'h00000647: inst = 32'h13058550;
30'h00000648: inst = 32'h23201500;
30'h00000649: inst = 32'hb7102121;
30'h0000064a: inst = 32'h938070c3;
30'h0000064b: inst = 32'h3705ff3f;
30'h0000064c: inst = 32'h1305c550;
30'h0000064d: inst = 32'h23201500;
30'h0000064e: inst = 32'hb7300500;
30'h0000064f: inst = 32'h938030b0;
30'h00000650: inst = 32'h3705ff3f;
30'h00000651: inst = 32'h13050551;
30'h00000652: inst = 32'h23201500;
30'h00000653: inst = 32'hb7108b11;
30'h00000654: inst = 32'h93803066;
30'h00000655: inst = 32'h3705ff3f;
30'h00000656: inst = 32'h13054551;
30'h00000657: inst = 32'h23201500;
30'h00000658: inst = 32'hb710c006;
30'h00000659: inst = 32'h938030f9;
30'h0000065a: inst = 32'h3705ff3f;
30'h0000065b: inst = 32'h13058551;
30'h0000065c: inst = 32'h23201500;
30'h0000065d: inst = 32'hb7801300;
30'h0000065e: inst = 32'h93803039;
30'h0000065f: inst = 32'h3705ff3f;
30'h00000660: inst = 32'h1305c551;
30'h00000661: inst = 32'h23201500;
30'h00000662: inst = 32'hb7102143;
30'h00000663: inst = 32'h938070d3;
30'h00000664: inst = 32'h3705ff3f;
30'h00000665: inst = 32'h13050552;
30'h00000666: inst = 32'h23201500;
30'h00000667: inst = 32'hb7600d01;
30'h00000668: inst = 32'h938030d1;
30'h00000669: inst = 32'h3705ff3f;
30'h0000066a: inst = 32'h13054552;
30'h0000066b: inst = 32'h23201500;
30'h0000066c: inst = 32'hb7106587;
30'h0000066d: inst = 32'h938070a3;
30'h0000066e: inst = 32'h3705ff3f;
30'h0000066f: inst = 32'h13058552;
30'h00000670: inst = 32'h23201500;
30'h00000671: inst = 32'hb7104d01;
30'h00000672: inst = 32'h9380309b;
30'h00000673: inst = 32'h3705ff3f;
30'h00000674: inst = 32'h1305c552;
30'h00000675: inst = 32'h23201500;
30'h00000676: inst = 32'hb7203501;
30'h00000677: inst = 32'h93803022;
30'h00000678: inst = 32'h3705ff3f;
30'h00000679: inst = 32'h13050553;
30'h0000067a: inst = 32'h23201500;
30'h0000067b: inst = 32'hb7304500;
30'h0000067c: inst = 32'h938030b0;
30'h0000067d: inst = 32'h3705ff3f;
30'h0000067e: inst = 32'h13054553;
30'h0000067f: inst = 32'h23201500;
30'h00000680: inst = 32'hb790690f;
30'h00000681: inst = 32'h93803046;
30'h00000682: inst = 32'h3705ff3f;
30'h00000683: inst = 32'h13058553;
30'h00000684: inst = 32'h23201500;
30'h00000685: inst = 32'hb710f006;
30'h00000686: inst = 32'h938030f9;
30'h00000687: inst = 32'h3705ff3f;
30'h00000688: inst = 32'h1305c553;
30'h00000689: inst = 32'h23201500;
30'h0000068a: inst = 32'hb7801300;
30'h0000068b: inst = 32'h93803039;
30'h0000068c: inst = 32'h3705ff3f;
30'h0000068d: inst = 32'h13050554;
30'h0000068e: inst = 32'h23201500;
30'h0000068f: inst = 32'hb7000010;
30'h00000690: inst = 32'h93807053;
30'h00000691: inst = 32'h3705ff3f;
30'h00000692: inst = 32'h13054554;
30'h00000693: inst = 32'h23201500;
30'h00000694: inst = 32'hb7102143;
30'h00000695: inst = 32'h938070d3;
30'h00000696: inst = 32'h3705ff3f;
30'h00000697: inst = 32'h13058554;
30'h00000698: inst = 32'h23201500;
30'h00000699: inst = 32'hb7600d01;
30'h0000069a: inst = 32'h938030d1;
30'h0000069b: inst = 32'h3705ff3f;
30'h0000069c: inst = 32'h1305c554;
30'h0000069d: inst = 32'h23201500;
30'h0000069e: inst = 32'hb7106587;
30'h0000069f: inst = 32'h938070a3;
30'h000006a0: inst = 32'h3705ff3f;
30'h000006a1: inst = 32'h13050555;
30'h000006a2: inst = 32'h23201500;
30'h000006a3: inst = 32'hb7104d01;
30'h000006a4: inst = 32'h9380309b;
30'h000006a5: inst = 32'h3705ff3f;
30'h000006a6: inst = 32'h13054555;
30'h000006a7: inst = 32'h23201500;
30'h000006a8: inst = 32'hb7203501;
30'h000006a9: inst = 32'h93803002;
30'h000006aa: inst = 32'h3705ff3f;
30'h000006ab: inst = 32'h13058555;
30'h000006ac: inst = 32'h23201500;
30'h000006ad: inst = 32'hb7103412;
30'h000006ae: inst = 32'h938070d3;
30'h000006af: inst = 32'h3705ff3f;
30'h000006b0: inst = 32'h1305c555;
30'h000006b1: inst = 32'h23201500;
30'h000006b2: inst = 32'hb7600d01;
30'h000006b3: inst = 32'h938030d1;
30'h000006b4: inst = 32'h3705ff3f;
30'h000006b5: inst = 32'h13050556;
30'h000006b6: inst = 32'h23201500;
30'h000006b7: inst = 32'hb710a501;
30'h000006b8: inst = 32'h93803002;
30'h000006b9: inst = 32'h3705ff3f;
30'h000006ba: inst = 32'h13054556;
30'h000006bb: inst = 32'h23201500;
30'h000006bc: inst = 32'hb7300500;
30'h000006bd: inst = 32'h938030b0;
30'h000006be: inst = 32'h3705ff3f;
30'h000006bf: inst = 32'h13058556;
30'h000006c0: inst = 32'h23201500;
30'h000006c1: inst = 32'hb7103412;
30'h000006c2: inst = 32'h938070d3;
30'h000006c3: inst = 32'h3705ff3f;
30'h000006c4: inst = 32'h1305c556;
30'h000006c5: inst = 32'h23201500;
30'h000006c6: inst = 32'hb7600d01;
30'h000006c7: inst = 32'h938030d1;
30'h000006c8: inst = 32'h3705ff3f;
30'h000006c9: inst = 32'h13050557;
30'h000006ca: inst = 32'h23201500;
30'h000006cb: inst = 32'hb7106587;
30'h000006cc: inst = 32'h938070a3;
30'h000006cd: inst = 32'h3705ff3f;
30'h000006ce: inst = 32'h13054557;
30'h000006cf: inst = 32'h23201500;
30'h000006d0: inst = 32'hb7104d01;
30'h000006d1: inst = 32'h938030c3;
30'h000006d2: inst = 32'h3705ff3f;
30'h000006d3: inst = 32'h13058557;
30'h000006d4: inst = 32'h23201500;
30'h000006d5: inst = 32'hb7108b0b;
30'h000006d6: inst = 32'h93803026;
30'h000006d7: inst = 32'h3705ff3f;
30'h000006d8: inst = 32'h1305c557;
30'h000006d9: inst = 32'h23201500;
30'h000006da: inst = 32'hb7102143;
30'h000006db: inst = 32'h938070d3;
30'h000006dc: inst = 32'h3705ff3f;
30'h000006dd: inst = 32'h13050558;
30'h000006de: inst = 32'h23201500;
30'h000006df: inst = 32'hb7600d01;
30'h000006e0: inst = 32'h938030d1;
30'h000006e1: inst = 32'h3705ff3f;
30'h000006e2: inst = 32'h13054558;
30'h000006e3: inst = 32'h23201500;
30'h000006e4: inst = 32'hb710a501;
30'h000006e5: inst = 32'h93803012;
30'h000006e6: inst = 32'h3705ff3f;
30'h000006e7: inst = 32'h13058558;
30'h000006e8: inst = 32'h23201500;
30'h000006e9: inst = 32'hb7300500;
30'h000006ea: inst = 32'h938030b0;
30'h000006eb: inst = 32'h3705ff3f;
30'h000006ec: inst = 32'h1305c558;
30'h000006ed: inst = 32'h23201500;
30'h000006ee: inst = 32'hb7103412;
30'h000006ef: inst = 32'h938070cb;
30'h000006f0: inst = 32'h3705ff3f;
30'h000006f1: inst = 32'h13050559;
30'h000006f2: inst = 32'h23201500;
30'h000006f3: inst = 32'hb7e00c01;
30'h000006f4: inst = 32'h938030c9;
30'h000006f5: inst = 32'h3705ff3f;
30'h000006f6: inst = 32'h13054559;
30'h000006f7: inst = 32'h23201500;
30'h000006f8: inst = 32'hb7102143;
30'h000006f9: inst = 32'h938070a3;
30'h000006fa: inst = 32'h3705ff3f;
30'h000006fb: inst = 32'h13058559;
30'h000006fc: inst = 32'h23201500;
30'h000006fd: inst = 32'hb7904c01;
30'h000006fe: inst = 32'h938030c3;
30'h000006ff: inst = 32'h3705ff3f;
30'h00000700: inst = 32'h1305c559;
30'h00000701: inst = 32'h23201500;
30'h00000702: inst = 32'hb7108b09;
30'h00000703: inst = 32'h93803006;
30'h00000704: inst = 32'h3705ff3f;
30'h00000705: inst = 32'h1305055a;
30'h00000706: inst = 32'h23201500;
30'h00000707: inst = 32'hb7100007;
30'h00000708: inst = 32'h938030f9;
30'h00000709: inst = 32'h3705ff3f;
30'h0000070a: inst = 32'h1305455a;
30'h0000070b: inst = 32'h23201500;
30'h0000070c: inst = 32'hb7801300;
30'h0000070d: inst = 32'h93803039;
30'h0000070e: inst = 32'h3705ff3f;
30'h0000070f: inst = 32'h1305855a;
30'h00000710: inst = 32'h23201500;
30'h00000711: inst = 32'hb7000010;
30'h00000712: inst = 32'h93807053;
30'h00000713: inst = 32'h3705ff3f;
30'h00000714: inst = 32'h1305c55a;
30'h00000715: inst = 32'h23201500;
30'h00000716: inst = 32'hb7004500;
30'h00000717: inst = 32'h93803059;
30'h00000718: inst = 32'h3705ff3f;
30'h00000719: inst = 32'h1305055b;
30'h0000071a: inst = 32'h23201500;
30'h0000071b: inst = 32'hb7105000;
30'h0000071c: inst = 32'h938030d1;
30'h0000071d: inst = 32'h3705ff3f;
30'h0000071e: inst = 32'h1305455b;
30'h0000071f: inst = 32'h23201500;
30'h00000720: inst = 32'hb7b0a5ff;
30'h00000721: inst = 32'h938030e2;
30'h00000722: inst = 32'h3705ff3f;
30'h00000723: inst = 32'h1305855b;
30'h00000724: inst = 32'h23201500;
30'h00000725: inst = 32'hb7200500;
30'h00000726: inst = 32'h93803028;
30'h00000727: inst = 32'h3705ff3f;
30'h00000728: inst = 32'h1305c55b;
30'h00000729: inst = 32'h23201500;
30'h0000072a: inst = 32'hb790a207;
30'h0000072b: inst = 32'h93803006;
30'h0000072c: inst = 32'h3705ff3f;
30'h0000072d: inst = 32'h1305055c;
30'h0000072e: inst = 32'h23201500;
30'h0000072f: inst = 32'hb7101007;
30'h00000730: inst = 32'h938030f9;
30'h00000731: inst = 32'h3705ff3f;
30'h00000732: inst = 32'h1305455c;
30'h00000733: inst = 32'h23201500;
30'h00000734: inst = 32'hb7801300;
30'h00000735: inst = 32'h93803039;
30'h00000736: inst = 32'h3705ff3f;
30'h00000737: inst = 32'h1305855c;
30'h00000738: inst = 32'h23201500;
30'h00000739: inst = 32'hb700c000;
30'h0000073a: inst = 32'h9380f00e;
30'h0000073b: inst = 32'h3705ff3f;
30'h0000073c: inst = 32'h1305c55c;
30'h0000073d: inst = 32'h23201500;
30'h0000073e: inst = 32'hb7a00500;
30'h0000073f: inst = 32'h93803040;
30'h00000740: inst = 32'h3705ff3f;
30'h00000741: inst = 32'h1305055d;
30'h00000742: inst = 32'h23201500;
30'h00000743: inst = 32'hb7106404;
30'h00000744: inst = 32'h93803066;
30'h00000745: inst = 32'h3705ff3f;
30'h00000746: inst = 32'h1305455d;
30'h00000747: inst = 32'h23201500;
30'h00000748: inst = 32'hb7006000;
30'h00000749: inst = 32'h93803031;
30'h0000074a: inst = 32'h3705ff3f;
30'h0000074b: inst = 32'h1305855d;
30'h0000074c: inst = 32'h23201500;
30'h0000074d: inst = 32'hb7000010;
30'h0000074e: inst = 32'h9380705b;
30'h0000074f: inst = 32'h3705ff3f;
30'h00000750: inst = 32'h1305c55d;
30'h00000751: inst = 32'h23201500;
30'h00000752: inst = 32'hb7000040;
30'h00000753: inst = 32'h93803051;
30'h00000754: inst = 32'h3705ff3f;
30'h00000755: inst = 32'h1305055e;
30'h00000756: inst = 32'h23201500;
30'h00000757: inst = 32'hb7108500;
30'h00000758: inst = 32'h93803051;
30'h00000759: inst = 32'h3705ff3f;
30'h0000075a: inst = 32'h1305455e;
30'h0000075b: inst = 32'h23201500;
30'h0000075c: inst = 32'hb700b500;
30'h0000075d: inst = 32'h9380305b;
30'h0000075e: inst = 32'h3705ff3f;
30'h0000075f: inst = 32'h1305855e;
30'h00000760: inst = 32'h23201500;
30'h00000761: inst = 32'hb7a06500;
30'h00000762: inst = 32'h93803002;
30'h00000763: inst = 32'h3705ff3f;
30'h00000764: inst = 32'h1305c55e;
30'h00000765: inst = 32'h23201500;
30'h00000766: inst = 32'hb7800000;
30'h00000767: inst = 32'h9380700e;
30'h00000768: inst = 32'h3705ff3f;
30'h00000769: inst = 32'h1305055f;
30'h0000076a: inst = 32'h23201500;
30'h0000076b: inst = 32'hb7102007;
30'h0000076c: inst = 32'h938030f9;
30'h0000076d: inst = 32'h3705ff3f;
30'h0000076e: inst = 32'h1305455f;
30'h0000076f: inst = 32'h23201500;
30'h00000770: inst = 32'hb7801300;
30'h00000771: inst = 32'h93803039;
30'h00000772: inst = 32'h3705ff3f;
30'h00000773: inst = 32'h1305855f;
30'h00000774: inst = 32'h23201500;
30'h00000775: inst = 32'hb7002000;
30'h00000776: inst = 32'h93803011;
30'h00000777: inst = 32'h3705ff3f;
30'h00000778: inst = 32'h1305c55f;
30'h00000779: inst = 32'h23201500;
30'h0000077a: inst = 32'hb7100000;
30'h0000077b: inst = 32'h938030a3;
30'h0000077c: inst = 32'h3705ff3f;
30'h0000077d: inst = 32'h13050560;
30'h0000077e: inst = 32'h23201500;
30'h0000077f: inst = 32'h93003046;
30'h00000780: inst = 32'h3705ff3f;
30'h00000781: inst = 32'h13054560;
30'h00000782: inst = 32'h23201500;
30'h00000783: inst = 32'hb710aa00;
30'h00000784: inst = 32'h938030a1;
30'h00000785: inst = 32'h3705ff3f;
30'h00000786: inst = 32'h13058560;
30'h00000787: inst = 32'h23201500;
30'h00000788: inst = 32'h93003003;
30'h00000789: inst = 32'h3705ff3f;
30'h0000078a: inst = 32'h1305c560;
30'h0000078b: inst = 32'h23201500;
30'h0000078c: inst = 32'h93003003;
30'h0000078d: inst = 32'h3705ff3f;
30'h0000078e: inst = 32'h13050561;
30'h0000078f: inst = 32'h23201500;
30'h00000790: inst = 32'hb7102a00;
30'h00000791: inst = 32'h938030a1;
30'h00000792: inst = 32'h3705ff3f;
30'h00000793: inst = 32'h13054561;
30'h00000794: inst = 32'h23201500;
30'h00000795: inst = 32'hb7104101;
30'h00000796: inst = 32'h93803046;
30'h00000797: inst = 32'h3705ff3f;
30'h00000798: inst = 32'h13058561;
30'h00000799: inst = 32'h23201500;
30'h0000079a: inst = 32'hb700c00e;
30'h0000079b: inst = 32'h9380f006;
30'h0000079c: inst = 32'h3705ff3f;
30'h0000079d: inst = 32'h1305c561;
30'h0000079e: inst = 32'h23201500;
30'h0000079f: inst = 32'hb7006004;
30'h000007a0: inst = 32'h93803021;
30'h000007a1: inst = 32'h3705ff3f;
30'h000007a2: inst = 32'h13050562;
30'h000007a3: inst = 32'h23201500;
30'h000007a4: inst = 32'hb7008017;
30'h000007a5: inst = 32'h9380f00e;
30'h000007a6: inst = 32'h3705ff3f;
30'h000007a7: inst = 32'h13054562;
30'h000007a8: inst = 32'h23201500;
30'h000007a9: inst = 32'hb7001004;
30'h000007aa: inst = 32'h93803021;
30'h000007ab: inst = 32'h3705ff3f;
30'h000007ac: inst = 32'h13058562;
30'h000007ad: inst = 32'h23201500;
30'h000007ae: inst = 32'hb7000017;
30'h000007af: inst = 32'h9380f00e;
30'h000007b0: inst = 32'h3705ff3f;
30'h000007b1: inst = 32'h1305c562;
30'h000007b2: inst = 32'h23201500;
30'h000007b3: inst = 32'hb7009004;
30'h000007b4: inst = 32'h93803021;
30'h000007b5: inst = 32'h3705ff3f;
30'h000007b6: inst = 32'h13050563;
30'h000007b7: inst = 32'h23201500;
30'h000007b8: inst = 32'hb7008016;
30'h000007b9: inst = 32'h9380f00e;
30'h000007ba: inst = 32'h3705ff3f;
30'h000007bb: inst = 32'h13054563;
30'h000007bc: inst = 32'h23201500;
30'h000007bd: inst = 32'hb700c004;
30'h000007be: inst = 32'h93803021;
30'h000007bf: inst = 32'h3705ff3f;
30'h000007c0: inst = 32'h13058563;
30'h000007c1: inst = 32'h23201500;
30'h000007c2: inst = 32'hb7000016;
30'h000007c3: inst = 32'h9380f00e;
30'h000007c4: inst = 32'h3705ff3f;
30'h000007c5: inst = 32'h1305c563;
30'h000007c6: inst = 32'h23201500;
30'h000007c7: inst = 32'hb7006004;
30'h000007c8: inst = 32'h93803021;
30'h000007c9: inst = 32'h3705ff3f;
30'h000007ca: inst = 32'h13050564;
30'h000007cb: inst = 32'h23201500;
30'h000007cc: inst = 32'hb7008015;
30'h000007cd: inst = 32'h9380f00e;
30'h000007ce: inst = 32'h3705ff3f;
30'h000007cf: inst = 32'h13054564;
30'h000007d0: inst = 32'h23201500;
30'h000007d1: inst = 32'hb7001004;
30'h000007d2: inst = 32'h93803021;
30'h000007d3: inst = 32'h3705ff3f;
30'h000007d4: inst = 32'h13058564;
30'h000007d5: inst = 32'h23201500;
30'h000007d6: inst = 32'hb7000015;
30'h000007d7: inst = 32'h9380f00e;
30'h000007d8: inst = 32'h3705ff3f;
30'h000007d9: inst = 32'h1305c564;
30'h000007da: inst = 32'h23201500;
30'h000007db: inst = 32'hb7009004;
30'h000007dc: inst = 32'h93803021;
30'h000007dd: inst = 32'h3705ff3f;
30'h000007de: inst = 32'h13050565;
30'h000007df: inst = 32'h23201500;
30'h000007e0: inst = 32'hb7008014;
30'h000007e1: inst = 32'h9380f00e;
30'h000007e2: inst = 32'h3705ff3f;
30'h000007e3: inst = 32'h13054565;
30'h000007e4: inst = 32'h23201500;
30'h000007e5: inst = 32'hb700c004;
30'h000007e6: inst = 32'h93803021;
30'h000007e7: inst = 32'h3705ff3f;
30'h000007e8: inst = 32'h13058565;
30'h000007e9: inst = 32'h23201500;
30'h000007ea: inst = 32'hb7000014;
30'h000007eb: inst = 32'h9380f00e;
30'h000007ec: inst = 32'h3705ff3f;
30'h000007ed: inst = 32'h1305c565;
30'h000007ee: inst = 32'h23201500;
30'h000007ef: inst = 32'hb7006004;
30'h000007f0: inst = 32'h93803021;
30'h000007f1: inst = 32'h3705ff3f;
30'h000007f2: inst = 32'h13050566;
30'h000007f3: inst = 32'h23201500;
30'h000007f4: inst = 32'hb7008013;
30'h000007f5: inst = 32'h9380f00e;
30'h000007f6: inst = 32'h3705ff3f;
30'h000007f7: inst = 32'h13054566;
30'h000007f8: inst = 32'h23201500;
30'h000007f9: inst = 32'hb7001004;
30'h000007fa: inst = 32'h93803021;
30'h000007fb: inst = 32'h3705ff3f;
30'h000007fc: inst = 32'h13058566;
30'h000007fd: inst = 32'h23201500;
30'h000007fe: inst = 32'hb7000013;
30'h000007ff: inst = 32'h9380f00e;
30'h00000800: inst = 32'h3705ff3f;
30'h00000801: inst = 32'h1305c566;
30'h00000802: inst = 32'h23201500;
30'h00000803: inst = 32'hb7009004;
30'h00000804: inst = 32'h93803021;
30'h00000805: inst = 32'h3705ff3f;
30'h00000806: inst = 32'h13050567;
30'h00000807: inst = 32'h23201500;
30'h00000808: inst = 32'hb7008012;
30'h00000809: inst = 32'h9380f00e;
30'h0000080a: inst = 32'h3705ff3f;
30'h0000080b: inst = 32'h13054567;
30'h0000080c: inst = 32'h23201500;
30'h0000080d: inst = 32'hb700c004;
30'h0000080e: inst = 32'h93803021;
30'h0000080f: inst = 32'h3705ff3f;
30'h00000810: inst = 32'h13058567;
30'h00000811: inst = 32'h23201500;
30'h00000812: inst = 32'hb7000012;
30'h00000813: inst = 32'h9380f00e;
30'h00000814: inst = 32'h3705ff3f;
30'h00000815: inst = 32'h1305c567;
30'h00000816: inst = 32'h23201500;
30'h00000817: inst = 32'hb7006004;
30'h00000818: inst = 32'h93803021;
30'h00000819: inst = 32'h3705ff3f;
30'h0000081a: inst = 32'h13050568;
30'h0000081b: inst = 32'h23201500;
30'h0000081c: inst = 32'hb7008011;
30'h0000081d: inst = 32'h9380f00e;
30'h0000081e: inst = 32'h3705ff3f;
30'h0000081f: inst = 32'h13054568;
30'h00000820: inst = 32'h23201500;
30'h00000821: inst = 32'hb7001004;
30'h00000822: inst = 32'h93803021;
30'h00000823: inst = 32'h3705ff3f;
30'h00000824: inst = 32'h13058568;
30'h00000825: inst = 32'h23201500;
30'h00000826: inst = 32'hb7000011;
30'h00000827: inst = 32'h9380f00e;
30'h00000828: inst = 32'h3705ff3f;
30'h00000829: inst = 32'h1305c568;
30'h0000082a: inst = 32'h23201500;
30'h0000082b: inst = 32'hb7009004;
30'h0000082c: inst = 32'h93803021;
30'h0000082d: inst = 32'h3705ff3f;
30'h0000082e: inst = 32'h13050569;
30'h0000082f: inst = 32'h23201500;
30'h00000830: inst = 32'hb7008010;
30'h00000831: inst = 32'h9380f00e;
30'h00000832: inst = 32'h3705ff3f;
30'h00000833: inst = 32'h13054569;
30'h00000834: inst = 32'h23201500;
30'h00000835: inst = 32'hb700c004;
30'h00000836: inst = 32'h93803021;
30'h00000837: inst = 32'h3705ff3f;
30'h00000838: inst = 32'h13058569;
30'h00000839: inst = 32'h23201500;
30'h0000083a: inst = 32'hb7000010;
30'h0000083b: inst = 32'h9380f00e;
30'h0000083c: inst = 32'h3705ff3f;
30'h0000083d: inst = 32'h1305c569;
30'h0000083e: inst = 32'h23201500;
30'h0000083f: inst = 32'hb700a003;
30'h00000840: inst = 32'h93803021;
30'h00000841: inst = 32'h3705ff3f;
30'h00000842: inst = 32'h1305056a;
30'h00000843: inst = 32'h23201500;
30'h00000844: inst = 32'hb700800f;
30'h00000845: inst = 32'h9380f00e;
30'h00000846: inst = 32'h3705ff3f;
30'h00000847: inst = 32'h1305456a;
30'h00000848: inst = 32'h23201500;
30'h00000849: inst = 32'hb7000002;
30'h0000084a: inst = 32'h93803021;
30'h0000084b: inst = 32'h3705ff3f;
30'h0000084c: inst = 32'h1305856a;
30'h0000084d: inst = 32'h23201500;
30'h0000084e: inst = 32'hb700000f;
30'h0000084f: inst = 32'h9380f00e;
30'h00000850: inst = 32'h3705ff3f;
30'h00000851: inst = 32'h1305c56a;
30'h00000852: inst = 32'h23201500;
30'h00000853: inst = 32'hb700f001;
30'h00000854: inst = 32'h93803023;
30'h00000855: inst = 32'h3705ff3f;
30'h00000856: inst = 32'h1305056b;
30'h00000857: inst = 32'h23201500;
30'h00000858: inst = 32'hb700800e;
30'h00000859: inst = 32'h9380f00e;
30'h0000085a: inst = 32'h3705ff3f;
30'h0000085b: inst = 32'h1305456b;
30'h0000085c: inst = 32'h23201500;
30'h0000085d: inst = 32'hb700a000;
30'h0000085e: inst = 32'h93803021;
30'h0000085f: inst = 32'h3705ff3f;
30'h00000860: inst = 32'h1305856b;
30'h00000861: inst = 32'h23201500;
30'h00000862: inst = 32'hb700000e;
30'h00000863: inst = 32'h9380f00e;
30'h00000864: inst = 32'h3705ff3f;
30'h00000865: inst = 32'h1305c56b;
30'h00000866: inst = 32'h23201500;
30'h00000867: inst = 32'hb700400d;
30'h00000868: inst = 32'h9380f006;
30'h00000869: inst = 32'h3705ff3f;
30'h0000086a: inst = 32'h1305056c;
30'h0000086b: inst = 32'h23201500;
30'h0000086c: inst = 32'hb7006004;
30'h0000086d: inst = 32'h93803021;
30'h0000086e: inst = 32'h3705ff3f;
30'h0000086f: inst = 32'h1305456c;
30'h00000870: inst = 32'h23201500;
30'h00000871: inst = 32'hb700400d;
30'h00000872: inst = 32'h9380f00e;
30'h00000873: inst = 32'h3705ff3f;
30'h00000874: inst = 32'h1305856c;
30'h00000875: inst = 32'h23201500;
30'h00000876: inst = 32'hb700c004;
30'h00000877: inst = 32'h93803021;
30'h00000878: inst = 32'h3705ff3f;
30'h00000879: inst = 32'h1305c56c;
30'h0000087a: inst = 32'h23201500;
30'h0000087b: inst = 32'hb700c00c;
30'h0000087c: inst = 32'h9380f00e;
30'h0000087d: inst = 32'h3705ff3f;
30'h0000087e: inst = 32'h1305056d;
30'h0000087f: inst = 32'h23201500;
30'h00000880: inst = 32'hb7001004;
30'h00000881: inst = 32'h93803021;
30'h00000882: inst = 32'h3705ff3f;
30'h00000883: inst = 32'h1305456d;
30'h00000884: inst = 32'h23201500;
30'h00000885: inst = 32'hb700400c;
30'h00000886: inst = 32'h9380f00e;
30'h00000887: inst = 32'h3705ff3f;
30'h00000888: inst = 32'h1305856d;
30'h00000889: inst = 32'h23201500;
30'h0000088a: inst = 32'hb7007004;
30'h0000088b: inst = 32'h93803021;
30'h0000088c: inst = 32'h3705ff3f;
30'h0000088d: inst = 32'h1305c56d;
30'h0000088e: inst = 32'h23201500;
30'h0000088f: inst = 32'hb700c00b;
30'h00000890: inst = 32'h9380f00e;
30'h00000891: inst = 32'h3705ff3f;
30'h00000892: inst = 32'h1305056e;
30'h00000893: inst = 32'h23201500;
30'h00000894: inst = 32'hb700a003;
30'h00000895: inst = 32'h93803021;
30'h00000896: inst = 32'h3705ff3f;
30'h00000897: inst = 32'h1305456e;
30'h00000898: inst = 32'h23201500;
30'h00000899: inst = 32'hb700400b;
30'h0000089a: inst = 32'h9380f00e;
30'h0000089b: inst = 32'h3705ff3f;
30'h0000089c: inst = 32'h1305856e;
30'h0000089d: inst = 32'h23201500;
30'h0000089e: inst = 32'hb7000002;
30'h0000089f: inst = 32'h93803021;
30'h000008a0: inst = 32'h3705ff3f;
30'h000008a1: inst = 32'h1305c56e;
30'h000008a2: inst = 32'h23201500;
30'h000008a3: inst = 32'hb700c00a;
30'h000008a4: inst = 32'h9380f00e;
30'h000008a5: inst = 32'h3705ff3f;
30'h000008a6: inst = 32'h1305056f;
30'h000008a7: inst = 32'h23201500;
30'h000008a8: inst = 32'hb700f001;
30'h000008a9: inst = 32'h93803023;
30'h000008aa: inst = 32'h3705ff3f;
30'h000008ab: inst = 32'h1305456f;
30'h000008ac: inst = 32'h23201500;
30'h000008ad: inst = 32'hb700400a;
30'h000008ae: inst = 32'h9380f00e;
30'h000008af: inst = 32'h3705ff3f;
30'h000008b0: inst = 32'h1305856f;
30'h000008b1: inst = 32'h23201500;
30'h000008b2: inst = 32'hb700a000;
30'h000008b3: inst = 32'h93803021;
30'h000008b4: inst = 32'h3705ff3f;
30'h000008b5: inst = 32'h1305c56f;
30'h000008b6: inst = 32'h23201500;
30'h000008b7: inst = 32'hb700c009;
30'h000008b8: inst = 32'h9380f00e;
30'h000008b9: inst = 32'h3705ff3f;
30'h000008ba: inst = 32'h13050570;
30'h000008bb: inst = 32'h23201500;
30'h000008bc: inst = 32'hb7000009;
30'h000008bd: inst = 32'h9380f006;
30'h000008be: inst = 32'h3705ff3f;
30'h000008bf: inst = 32'h13054570;
30'h000008c0: inst = 32'h23201500;
30'h000008c1: inst = 32'hb7000005;
30'h000008c2: inst = 32'h93803021;
30'h000008c3: inst = 32'h3705ff3f;
30'h000008c4: inst = 32'h13058570;
30'h000008c5: inst = 32'h23201500;
30'h000008c6: inst = 32'hb7000009;
30'h000008c7: inst = 32'h9380f00e;
30'h000008c8: inst = 32'h3705ff3f;
30'h000008c9: inst = 32'h1305c570;
30'h000008ca: inst = 32'h23201500;
30'h000008cb: inst = 32'hb7001004;
30'h000008cc: inst = 32'h93803021;
30'h000008cd: inst = 32'h3705ff3f;
30'h000008ce: inst = 32'h13050571;
30'h000008cf: inst = 32'h23201500;
30'h000008d0: inst = 32'hb7008008;
30'h000008d1: inst = 32'h9380f00e;
30'h000008d2: inst = 32'h3705ff3f;
30'h000008d3: inst = 32'h13054571;
30'h000008d4: inst = 32'h23201500;
30'h000008d5: inst = 32'hb7003005;
30'h000008d6: inst = 32'h93803021;
30'h000008d7: inst = 32'h3705ff3f;
30'h000008d8: inst = 32'h13058571;
30'h000008d9: inst = 32'h23201500;
30'h000008da: inst = 32'hb7000008;
30'h000008db: inst = 32'h9380f00e;
30'h000008dc: inst = 32'h3705ff3f;
30'h000008dd: inst = 32'h1305c571;
30'h000008de: inst = 32'h23201500;
30'h000008df: inst = 32'hb7003005;
30'h000008e0: inst = 32'h93803021;
30'h000008e1: inst = 32'h3705ff3f;
30'h000008e2: inst = 32'h13050572;
30'h000008e3: inst = 32'h23201500;
30'h000008e4: inst = 32'hb7008007;
30'h000008e5: inst = 32'h9380f00e;
30'h000008e6: inst = 32'h3705ff3f;
30'h000008e7: inst = 32'h13054572;
30'h000008e8: inst = 32'h23201500;
30'h000008e9: inst = 32'hb7000005;
30'h000008ea: inst = 32'h93803021;
30'h000008eb: inst = 32'h3705ff3f;
30'h000008ec: inst = 32'h13058572;
30'h000008ed: inst = 32'h23201500;
30'h000008ee: inst = 32'hb7000007;
30'h000008ef: inst = 32'h9380f00e;
30'h000008f0: inst = 32'h3705ff3f;
30'h000008f1: inst = 32'h1305c572;
30'h000008f2: inst = 32'h23201500;
30'h000008f3: inst = 32'hb7001004;
30'h000008f4: inst = 32'h93803021;
30'h000008f5: inst = 32'h3705ff3f;
30'h000008f6: inst = 32'h13050573;
30'h000008f7: inst = 32'h23201500;
30'h000008f8: inst = 32'hb7008006;
30'h000008f9: inst = 32'h9380f00e;
30'h000008fa: inst = 32'h3705ff3f;
30'h000008fb: inst = 32'h13054573;
30'h000008fc: inst = 32'h23201500;
30'h000008fd: inst = 32'hb7003005;
30'h000008fe: inst = 32'h93803021;
30'h000008ff: inst = 32'h3705ff3f;
30'h00000900: inst = 32'h13058573;
30'h00000901: inst = 32'h23201500;
30'h00000902: inst = 32'hb7000006;
30'h00000903: inst = 32'h9380f00e;
30'h00000904: inst = 32'h3705ff3f;
30'h00000905: inst = 32'h1305c573;
30'h00000906: inst = 32'h23201500;
30'h00000907: inst = 32'hb7003005;
30'h00000908: inst = 32'h93803021;
30'h00000909: inst = 32'h3705ff3f;
30'h0000090a: inst = 32'h13050574;
30'h0000090b: inst = 32'h23201500;
30'h0000090c: inst = 32'hb7008005;
30'h0000090d: inst = 32'h9380f00e;
30'h0000090e: inst = 32'h3705ff3f;
30'h0000090f: inst = 32'h13054574;
30'h00000910: inst = 32'h23201500;
30'h00000911: inst = 32'hb7000005;
30'h00000912: inst = 32'h93803021;
30'h00000913: inst = 32'h3705ff3f;
30'h00000914: inst = 32'h13058574;
30'h00000915: inst = 32'h23201500;
30'h00000916: inst = 32'hb7000005;
30'h00000917: inst = 32'h9380f00e;
30'h00000918: inst = 32'h3705ff3f;
30'h00000919: inst = 32'h1305c574;
30'h0000091a: inst = 32'h23201500;
30'h0000091b: inst = 32'hb7001004;
30'h0000091c: inst = 32'h93803021;
30'h0000091d: inst = 32'h3705ff3f;
30'h0000091e: inst = 32'h13050575;
30'h0000091f: inst = 32'h23201500;
30'h00000920: inst = 32'hb7008004;
30'h00000921: inst = 32'h9380f00e;
30'h00000922: inst = 32'h3705ff3f;
30'h00000923: inst = 32'h13054575;
30'h00000924: inst = 32'h23201500;
30'h00000925: inst = 32'hb7003005;
30'h00000926: inst = 32'h93803021;
30'h00000927: inst = 32'h3705ff3f;
30'h00000928: inst = 32'h13058575;
30'h00000929: inst = 32'h23201500;
30'h0000092a: inst = 32'hb7000004;
30'h0000092b: inst = 32'h9380f00e;
30'h0000092c: inst = 32'h3705ff3f;
30'h0000092d: inst = 32'h1305c575;
30'h0000092e: inst = 32'h23201500;
30'h0000092f: inst = 32'hb7003005;
30'h00000930: inst = 32'h93803021;
30'h00000931: inst = 32'h3705ff3f;
30'h00000932: inst = 32'h13050576;
30'h00000933: inst = 32'h23201500;
30'h00000934: inst = 32'hb7008003;
30'h00000935: inst = 32'h9380f00e;
30'h00000936: inst = 32'h3705ff3f;
30'h00000937: inst = 32'h13054576;
30'h00000938: inst = 32'h23201500;
30'h00000939: inst = 32'hb7000005;
30'h0000093a: inst = 32'h93803021;
30'h0000093b: inst = 32'h3705ff3f;
30'h0000093c: inst = 32'h13058576;
30'h0000093d: inst = 32'h23201500;
30'h0000093e: inst = 32'hb7000003;
30'h0000093f: inst = 32'h9380f00e;
30'h00000940: inst = 32'h3705ff3f;
30'h00000941: inst = 32'h1305c576;
30'h00000942: inst = 32'h23201500;
30'h00000943: inst = 32'hb7001004;
30'h00000944: inst = 32'h93803021;
30'h00000945: inst = 32'h3705ff3f;
30'h00000946: inst = 32'h13050577;
30'h00000947: inst = 32'h23201500;
30'h00000948: inst = 32'hb7008002;
30'h00000949: inst = 32'h9380f00e;
30'h0000094a: inst = 32'h3705ff3f;
30'h0000094b: inst = 32'h13054577;
30'h0000094c: inst = 32'h23201500;
30'h0000094d: inst = 32'hb7003005;
30'h0000094e: inst = 32'h93803021;
30'h0000094f: inst = 32'h3705ff3f;
30'h00000950: inst = 32'h13058577;
30'h00000951: inst = 32'h23201500;
30'h00000952: inst = 32'hb7000002;
30'h00000953: inst = 32'h9380f00e;
30'h00000954: inst = 32'h3705ff3f;
30'h00000955: inst = 32'h1305c577;
30'h00000956: inst = 32'h23201500;
30'h00000957: inst = 32'hb7003005;
30'h00000958: inst = 32'h93803021;
30'h00000959: inst = 32'h3705ff3f;
30'h0000095a: inst = 32'h13050578;
30'h0000095b: inst = 32'h23201500;
30'h0000095c: inst = 32'hb7008001;
30'h0000095d: inst = 32'h9380f00e;
30'h0000095e: inst = 32'h3705ff3f;
30'h0000095f: inst = 32'h13054578;
30'h00000960: inst = 32'h23201500;
30'h00000961: inst = 32'hb700a000;
30'h00000962: inst = 32'h93803021;
30'h00000963: inst = 32'h3705ff3f;
30'h00000964: inst = 32'h13058578;
30'h00000965: inst = 32'h23201500;
30'h00000966: inst = 32'hb7000001;
30'h00000967: inst = 32'h9380f00e;
30'h00000968: inst = 32'h3705ff3f;
30'h00000969: inst = 32'h1305c578;
30'h0000096a: inst = 32'h23201500;
30'h0000096b: inst = 32'hb7004000;
30'h0000096c: inst = 32'h9380f006;
30'h0000096d: inst = 32'h3705ff3f;
30'h0000096e: inst = 32'h13050579;
30'h0000096f: inst = 32'h23201500;
30'h00000970: inst = 32'hb7101000;
30'h00000971: inst = 32'h938030f1;
30'h00000972: inst = 32'h3705ff3f;
30'h00000973: inst = 32'h13054579;
30'h00000974: inst = 32'h23201500;
30'h00000975: inst = 32'hb7f0dfff;
30'h00000976: inst = 32'h9380f006;
30'h00000977: inst = 32'h3705ff3f;
30'h00000978: inst = 32'h13058579;
30'h00000979: inst = 32'h23201500;
30'h0000097a: inst = 32'hb7000080;
30'h0000097b: inst = 32'h93807013;
30'h0000097c: inst = 32'h3705ff3f;
30'h0000097d: inst = 32'h1305c579;
30'h0000097e: inst = 32'h23201500;
30'h0000097f: inst = 32'hb7200100;
30'h00000980: inst = 32'h93803018;
30'h00000981: inst = 32'h3705ff3f;
30'h00000982: inst = 32'h1305057a;
30'h00000983: inst = 32'h23201500;
30'h00000984: inst = 32'hb7f01100;
30'h00000985: inst = 32'h93803019;
30'h00000986: inst = 32'h3705ff3f;
30'h00000987: inst = 32'h1305457a;
30'h00000988: inst = 32'h23201500;
30'h00000989: inst = 32'hb79001fe;
30'h0000098a: inst = 32'h938030ae;
30'h0000098b: inst = 32'h3705ff3f;
30'h0000098c: inst = 32'h1305857a;
30'h0000098d: inst = 32'h23201500;
30'h0000098e: inst = 32'hb7204100;
30'h0000098f: inst = 32'h93803042;
30'h00000990: inst = 32'h3705ff3f;
30'h00000991: inst = 32'h1305c57a;
30'h00000992: inst = 32'h23201500;
30'h00000993: inst = 32'hb7800000;
30'h00000994: inst = 32'h93807006;
30'h00000995: inst = 32'h3705ff3f;
30'h00000996: inst = 32'h1305057b;
30'h00000997: inst = 32'h23201500;
30'h00000998: inst = 32'h3705ff1f;
30'h00000999: inst = 32'h67000500;
default:      inst = 32'h00000000;
endcase
end
endmodule
